    always @(dq_in[45]) dq_timing_check(45);