    always @(addr[1]) addr_timing_check(1);