    always @(posedge ck) begin
        audio_raddr_0 <= audio_raddr;
    end