    always @(dq_in[33]) dq_timing_check(33);