	 always @(*)
		if (control)
			c = b;
		else
			c = a;
		