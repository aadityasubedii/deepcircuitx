    always @(addr[0]) addr_timing_check(0);
