    always @(dm_in[14]) dm_timing_check(14);