  always@(posedge clk, posedge reset) begin
    if(reset) begin 
      Y     <= RSTVAL; 
      R[30] <= RSTVAL;
      R[29] <= RSTVAL;
      R[28] <= RSTVAL;
      R[27] <= RSTVAL;
      R[26] <= RSTVAL;
      R[25] <= RSTVAL;
      R[24] <= RSTVAL;
      R[23] <= RSTVAL;
      R[22] <= RSTVAL;
      R[21] <= RSTVAL;
      R[20] <= RSTVAL;
      R[19] <= RSTVAL;
      R[18] <= RSTVAL;
      R[17] <= RSTVAL;
      R[16] <= RSTVAL;
      R[15] <= RSTVAL;
      R[14] <= RSTVAL;
      R[13] <= RSTVAL;
      R[12] <= RSTVAL;
      R[11] <= RSTVAL;
      R[10] <= RSTVAL;
      R[9]  <= RSTVAL;
      R[8]  <= RSTVAL;
      R[7]  <= RSTVAL;
      R[6]  <= RSTVAL;
      R[5]  <= RSTVAL;
      R[4]  <= RSTVAL;
      R[3]  <= RSTVAL;
      R[2]  <= RSTVAL;
      R[1]  <= RSTVAL;
      R[0]  <= RSTVAL;
    end
    else begin 
      Y     <= R[30];
      R[30] <= R[29];
      R[29] <= R[28];
      R[28] <= R[27];
      R[27] <= R[26];
      R[26] <= R[25];
      R[25] <= R[24];
      R[24] <= R[23];
      R[23] <= R[22];
      R[22] <= R[21];
      R[21] <= R[20];
      R[20] <= R[19];
      R[19] <= R[18];
      R[18] <= R[17];
      R[17] <= R[16];
      R[16] <= R[15];
      R[15] <= R[14];
      R[14] <= R[13];
      R[13] <= R[12];
      R[12] <= R[11];
      R[11] <= R[10];
      R[10] <= R[9];
      R[9]  <= R[8];
      R[8]  <= R[7];
      R[7]  <= R[6];
      R[6]  <= R[5];
      R[5]  <= R[4];
      R[4]  <= R[3];
      R[3]  <= R[2];
      R[2]  <= R[1];
      R[1]  <= R[0];
      R[0]  <= X;
    end
  end