module lab7_soc_nios2_gen2_0_cpu_nios2_oci_compute_input_tm_cnt (
                                                                  
                                                                   atm_valid,
                                                                   dtm_valid,
                                                                   itm_valid,

                                                                  
                                                                   compute_input_tm_cnt
                                                                )
;