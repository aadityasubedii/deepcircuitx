module delay4k(
  input wire [3:0] index,
  
output reg [11:0] delay
);