    always @(posedge dqs_in[18]) dqs_neg_timing_check(18);