    always @(posedge clk) sync_1 <= sync_0;