module lab7_soc_nios2_gen2_0_cpu_nios2_oci_im (
                                                
                                                 clk,
                                                 jrst_n,
                                                 trc_ctrl,
                                                 tw,

                                                
                                                 tracemem_on,
                                                 tracemem_trcdata,
                                                 tracemem_tw,
                                                 trc_im_addr,
                                                 trc_wrap,
                                                 xbrk_wrap_traceoff
                                              )