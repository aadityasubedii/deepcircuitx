            always @(posedge ck) begin
                delay <= in;
            end