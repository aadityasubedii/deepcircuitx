    always @(dq_in[31]) dq_timing_check(31);