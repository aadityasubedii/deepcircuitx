



endmodule