	always @ (posedge CLOCK_50)
		if (load == 1'b1) d <= SW;