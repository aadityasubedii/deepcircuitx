`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:46:09 08/20/2022 
// Design Name: 
// Module Name:    IN_IIR 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ECHO(clk, DATA_IN, DATA_OUT);

input clk;
input[11:0] DATA_IN;
output reg[11:0] DATA_OUT;

//wire signed[11:0] DATA_IN;

reg signed[11:0] IN[40:0];

initial begin

DATA_OUT = 12'b000000000000;
IN[0] = 12'b000000000000;
IN[1] = 12'b000000000000;
IN[2] = 12'b000000000000;
IN[3] = 12'b000000000000;
IN[4] = 12'b000000000000;
IN[5] = 12'b000000000000;
IN[6] = 12'b000000000000;
IN[7] = 12'b000000000000;
IN[8] = 12'b000000000000;
IN[9] = 12'b000000000000;
IN[10] = 12'b000000000000;
IN[11] = 12'b000000000000;
IN[12] = 12'b000000000000;
IN[13] = 12'b000000000000;
IN[14] = 12'b000000000000;
IN[15] = 12'b000000000000;
IN[16] = 12'b000000000000;
IN[17] = 12'b000000000000;
IN[18] = 12'b000000000000;
IN[19] = 12'b000000000000;
IN[20] = 12'b000000000000;
IN[21] = 12'b000000000000;
IN[22] = 12'b000000000000;
IN[23] = 12'b000000000000;
IN[24] = 12'b000000000000;
IN[25] = 12'b000000000000;
IN[26] = 12'b000000000000;
IN[27] = 12'b000000000000;
IN[28] = 12'b000000000000;
IN[29] = 12'b000000000000;
IN[30] = 12'b000000000000;
IN[31] = 12'b000000000000;
IN[32] = 12'b000000000000;
IN[33] = 12'b000000000000;
IN[34] = 12'b000000000000;
IN[35] = 12'b000000000000;
IN[36] = 12'b000000000000;
IN[37] = 12'b000000000000;
IN[38] = 12'b000000000000;
IN[39] = 12'b000000000000;
IN[40] = 12'b000000000000;

end

always@(DATA_IN)
begin
    DATA_OUT = DATA_IN + (IN[40]>>2 + IN[40]>>1);
end

always@(posedge clk)
begin
	
		IN[0] <= DATA_IN;
		IN[1] <= IN[0];
		IN[2] <= IN[1];
		IN[3] <= IN[2];
		IN[4] <= IN[3];
		IN[5] <= IN[4];
		IN[6] <= IN[5];
		IN[7] <= IN[6];
		IN[8] <= IN[7];
		IN[9] <= IN[8];
		IN[10] <= IN[9];
		IN[11] <= IN[10];
		IN[12] <= IN[11];
		IN[13] <= IN[12];
		IN[14] <= IN[13];
		IN[15] <= IN[14];
		IN[16] <= IN[15];
		IN[17] <= IN[16];
		IN[18] <= IN[17];
		IN[19] <= IN[18];
		IN[20] <= IN[19];
		IN[21] <= IN[20];
        IN[22] <= IN[21];
        IN[23] <= IN[22];
        IN[24] <= IN[23];
        IN[25] <= IN[24];
        IN[26] <= IN[25];
        IN[27] <= IN[26];
        IN[28] <= IN[27];
        IN[29] <= IN[28];
        IN[30] <= IN[29];
        IN[31] <= IN[30];
        IN[32] <= IN[31];
        IN[33] <= IN[32];
        IN[34] <= IN[33];
        IN[35] <= IN[34];
        IN[36] <= IN[35];
        IN[37] <= IN[36];
        IN[38] <= IN[37];
        IN[39] <= IN[38];
        IN[40] <= IN[39];

end
endmodule
