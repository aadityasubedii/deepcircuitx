`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/25/2023 10:51:38 PM
// Design Name: 
// Module Name: add_sub
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module add_sub(
    input [3:0] A, B,
    input en,
    output [3:0] sdout,
    output cbout
    );
    
    wire [2:0]c;
    
    full_adder fa1(A[0], (B[0]^en), en, sdout[0], c[0]);
    full_adder fa2(A[1], (B[1]^en), c[0], sdout[1], c[1]);
    full_adder fa3(A[2], (B[2]^en), c[1], sdout[2], c[2]);
    full_adder fa4(A[3], (B[3]^en), c[2], sdout[3], cbout);
 
endmodule
