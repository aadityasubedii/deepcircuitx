    always @(ba     ) ba_in      <= #BUS_DELAY ba;