
//Verilog file of module maxAbsValueCir


`timescale 1 ns / 1ns

module maxAbsValueCir_net(w1,
w2,
w3,
out);
input [0:3]w1;
input [0:3]w2;
input [0:3]w3;
output [0:3]out;
wire
maxAbsValueCir_wire_1,
maxAbsValueCir_wire_2,
maxAbsValueCir_wire_3,
maxAbsValueCir_wire_4,
maxAbsValueCir_wire_5,
maxAbsValueCir_wire_6,
maxAbsValueCir_wire_7,
maxAbsValueCir_wire_8,
maxAbsValueCir_wire_9,
maxAbsValueCir_wire_10,
maxAbsValueCir_wire_11,
maxAbsValueCir_wire_12,
maxAbsValueCir_wire_13,
maxAbsValueCir_wire_14,
maxAbsValueCir_wire_15,
maxAbsValueCir_wire_16,
maxAbsValueCir_wire_17,
maxAbsValueCir_wire_18,
maxAbsValueCir_wire_19,
maxAbsValueCir_wire_20,
maxAbsValueCir_wire_21,
maxAbsValueCir_wire_22,
maxAbsValueCir_wire_23,
maxAbsValueCir_wire_24,
maxAbsValueCir_wire_25,
maxAbsValueCir_wire_26,
maxAbsValueCir_wire_27,
maxAbsValueCir_wire_28,
maxAbsValueCir_wire_29,
maxAbsValueCir_wire_30,
maxAbsValueCir_wire_31,
maxAbsValueCir_wire_32,
maxAbsValueCir_wire_33,
maxAbsValueCir_wire_34,
maxAbsValueCir_wire_35,
maxAbsValueCir_wire_36,
maxAbsValueCir_wire_37,
maxAbsValueCir_wire_38,
maxAbsValueCir_wire_39,
maxAbsValueCir_wire_40,
maxAbsValueCir_wire_41,
maxAbsValueCir_wire_42,
maxAbsValueCir_wire_43,
maxAbsValueCir_wire_44,
maxAbsValueCir_wire_45,
maxAbsValueCir_wire_46,
maxAbsValueCir_wire_47,
maxAbsValueCir_wire_48,
maxAbsValueCir_wire_49,
maxAbsValueCir_wire_50,
maxAbsValueCir_wire_51,
maxAbsValueCir_wire_52,
maxAbsValueCir_wire_53,
maxAbsValueCir_wire_54,
maxAbsValueCir_wire_55,
maxAbsValueCir_wire_56,
maxAbsValueCir_wire_57,
maxAbsValueCir_wire_58,
maxAbsValueCir_wire_59,
maxAbsValueCir_wire_60,
maxAbsValueCir_wire_61,
maxAbsValueCir_wire_62,
maxAbsValueCir_wire_63,
maxAbsValueCir_wire_64,
maxAbsValueCir_wire_65,
maxAbsValueCir_wire_66,
maxAbsValueCir_wire_67,
maxAbsValueCir_wire_68,
maxAbsValueCir_wire_69,
maxAbsValueCir_wire_70,
maxAbsValueCir_wire_71,
maxAbsValueCir_wire_72,
maxAbsValueCir_wire_73,
maxAbsValueCir_wire_74,
maxAbsValueCir_wire_75,
maxAbsValueCir_wire_76,
maxAbsValueCir_wire_77,
maxAbsValueCir_wire_78,
maxAbsValueCir_wire_79,
maxAbsValueCir_wire_80,
maxAbsValueCir_wire_81,
maxAbsValueCir_wire_82,
maxAbsValueCir_wire_83,
maxAbsValueCir_wire_84,
maxAbsValueCir_wire_85,
maxAbsValueCir_wire_86,
maxAbsValueCir_wire_87,
maxAbsValueCir_wire_88,
maxAbsValueCir_wire_89,
maxAbsValueCir_wire_90,
maxAbsValueCir_wire_91,
maxAbsValueCir_wire_92,
maxAbsValueCir_wire_93,
maxAbsValueCir_wire_94,
maxAbsValueCir_wire_95,
maxAbsValueCir_wire_96,
maxAbsValueCir_wire_97,
maxAbsValueCir_wire_98,
maxAbsValueCir_wire_99,
maxAbsValueCir_wire_100,
maxAbsValueCir_wire_101,
maxAbsValueCir_wire_102,
maxAbsValueCir_wire_103,
maxAbsValueCir_wire_104,
maxAbsValueCir_wire_105,
maxAbsValueCir_wire_106,
maxAbsValueCir_wire_107,
maxAbsValueCir_wire_108,
maxAbsValueCir_wire_109,
maxAbsValueCir_wire_110,
maxAbsValueCir_wire_111,
maxAbsValueCir_wire_112,
maxAbsValueCir_wire_113,
maxAbsValueCir_wire_114,
maxAbsValueCir_wire_115,
maxAbsValueCir_wire_116,
maxAbsValueCir_wire_117,
maxAbsValueCir_wire_118,
maxAbsValueCir_wire_119,
maxAbsValueCir_wire_120,
maxAbsValueCir_wire_121,
maxAbsValueCir_wire_122,
maxAbsValueCir_wire_123,
maxAbsValueCir_wire_124,
maxAbsValueCir_wire_125,
maxAbsValueCir_wire_126,
maxAbsValueCir_wire_127,
maxAbsValueCir_wire_128,
maxAbsValueCir_wire_129,
maxAbsValueCir_wire_130,
maxAbsValueCir_wire_131,
maxAbsValueCir_wire_132,
maxAbsValueCir_wire_133,
maxAbsValueCir_wire_134,
maxAbsValueCir_wire_135,
maxAbsValueCir_wire_7_0,
maxAbsValueCir_wire_7_1,
maxAbsValueCir_wire_7_2,
maxAbsValueCir_wire_25_0,
maxAbsValueCir_wire_25_1,
maxAbsValueCir_wire_25_2,
maxAbsValueCir_wire_14_0,
maxAbsValueCir_wire_14_1,
maxAbsValueCir_wire_5_0,
maxAbsValueCir_wire_5_1,
maxAbsValueCir_wire_23_0,
maxAbsValueCir_wire_23_1,
maxAbsValueCir_wire_57_0,
maxAbsValueCir_wire_57_1,
maxAbsValueCir_wire_57_2,
maxAbsValueCir_wire_57_3,
maxAbsValueCir_wire_57_4,
maxAbsValueCir_wire_57_5,
maxAbsValueCir_wire_57_6,
maxAbsValueCir_wire_57_7,
maxAbsValueCir_wire_85_0,
maxAbsValueCir_wire_85_1,
maxAbsValueCir_wire_85_2,
maxAbsValueCir_wire_85_3,
maxAbsValueCir_wire_85_4,
maxAbsValueCir_wire_85_5,
maxAbsValueCir_wire_85_6,
maxAbsValueCir_wire_85_7,
maxAbsValueCir_wire_59_0,
maxAbsValueCir_wire_59_1,
maxAbsValueCir_wire_59_2,
maxAbsValueCir_wire_59_3,
maxAbsValueCir_wire_58_0,
maxAbsValueCir_wire_58_1,
maxAbsValueCir_wire_58_2,
maxAbsValueCir_wire_58_3,
maxAbsValueCir_wire_34_0,
maxAbsValueCir_wire_34_1,
maxAbsValueCir_wire_34_2,
maxAbsValueCir_wire_34_3,
maxAbsValueCir_wire_34_4,
maxAbsValueCir_wire_34_5,
maxAbsValueCir_wire_53_0,
maxAbsValueCir_wire_53_1,
maxAbsValueCir_wire_44_0,
maxAbsValueCir_wire_44_1,
maxAbsValueCir_wire_81_0,
maxAbsValueCir_wire_81_1,
maxAbsValueCir_wire_72_0,
maxAbsValueCir_wire_72_1,
maxAbsValueCir_wire_11_0,
maxAbsValueCir_wire_11_1,
maxAbsValueCir_wire_11_2,
maxAbsValueCir_wire_11_3,
maxAbsValueCir_wire_11_4,
maxAbsValueCir_wire_12_0,
maxAbsValueCir_wire_12_1,
maxAbsValueCir_wire_12_2,
maxAbsValueCir_wire_12_3,
maxAbsValueCir_wire_15_0,
maxAbsValueCir_wire_15_1,
maxAbsValueCir_wire_15_2,
maxAbsValueCir_wire_15_3,
maxAbsValueCir_wire_18_0,
maxAbsValueCir_wire_18_1,
maxAbsValueCir_wire_18_2,
maxAbsValueCir_wire_18_3,
maxAbsValueCir_wire_18_4,
maxAbsValueCir_wire_18_5,
maxAbsValueCir_wire_18_6,
maxAbsValueCir_wire_2_0,
maxAbsValueCir_wire_2_1,
maxAbsValueCir_wire_2_2,
maxAbsValueCir_wire_2_3,
maxAbsValueCir_wire_3_0,
maxAbsValueCir_wire_3_1,
maxAbsValueCir_wire_3_2,
maxAbsValueCir_wire_3_3,
maxAbsValueCir_wire_6_0,
maxAbsValueCir_wire_6_1,
maxAbsValueCir_wire_6_2,
maxAbsValueCir_wire_6_3,
maxAbsValueCir_wire_9_0,
maxAbsValueCir_wire_9_1,
maxAbsValueCir_wire_9_2,
maxAbsValueCir_wire_9_3,
maxAbsValueCir_wire_9_4,
maxAbsValueCir_wire_9_5,
maxAbsValueCir_wire_9_6,
maxAbsValueCir_wire_9_7,
maxAbsValueCir_wire_9_8,
maxAbsValueCir_wire_20_0,
maxAbsValueCir_wire_20_1,
maxAbsValueCir_wire_20_2,
maxAbsValueCir_wire_20_3,
maxAbsValueCir_wire_21_0,
maxAbsValueCir_wire_21_1,
maxAbsValueCir_wire_21_2,
maxAbsValueCir_wire_21_3,
maxAbsValueCir_wire_24_0,
maxAbsValueCir_wire_24_1,
maxAbsValueCir_wire_24_2,
maxAbsValueCir_wire_24_3,
maxAbsValueCir_wire_27_0,
maxAbsValueCir_wire_27_1,
maxAbsValueCir_wire_27_2,
maxAbsValueCir_wire_27_3,
maxAbsValueCir_wire_27_4,
maxAbsValueCir_wire_27_5,
maxAbsValueCir_wire_27_6,
maxAbsValueCir_wire_27_7,
maxAbsValueCir_wire_27_8;

pin #(12) pin_0 ({w1[0], w1[1], w1[2], w1[3], w2[0], w2[1], w2[2], w2[3], w3[0], w3[1], w3[2], w3[3]}, {w1_0, w1_1, w1_2, w1_3, w2_0, w2_1, w2_2, w2_3, w3_0, w3_1, w3_2, w3_3});

pout #(1108) pout_0 ({out_0, out_1, out_2, out_3, out_4, out_5, out_6, out_7, out_8, out_9, out_10, out_11, out_12, out_13, out_14, out_15, out_16, out_17, out_18, out_19, out_20, out_21, out_22, out_23, out_24, out_25, out_26, out_27, out_28, out_29, out_30, out_31, out_32, out_33, out_34, out_35, out_36, out_37, out_38, out_39, out_40, out_41, out_42, out_43, out_44, out_45, out_46, out_47, out_48, out_49, out_50, out_51, out_52, out_53, out_54, out_55, out_56, out_57, out_58, out_59, out_60, out_61, out_62, out_63, out_64, out_65, out_66, out_67, out_68, out_69, out_70, out_71, out_72, out_73, out_74, out_75, out_76, out_77, out_78, out_79, out_80, out_81, out_82, out_83, out_84, out_85, out_86, out_87, out_88, out_89, out_90, out_91, out_92, out_93, out_94, out_95, out_96, out_97, out_98, out_99, out_100, out_101, out_102, out_103, out_104, out_105, out_106, out_107, out_108, out_109, out_110, out_111, out_112, out_113, out_114, out_115, out_116, out_117, out_118, out_119, out_120, out_121, out_122, out_123, out_124, out_125, out_126, out_127, out_128, out_129, out_130, out_131, out_132, out_133, out_134, out_135, out_136, out_137, out_138, out_139, out_140, out_141, out_142, out_143, out_144, out_145, out_146, out_147, out_148, out_149, out_150, out_151, out_152, out_153, out_154, out_155, out_156, out_157, out_158, out_159, out_160, out_161, out_162, out_163, out_164, out_165, out_166, out_167, out_168, out_169, out_170, out_171, out_172, out_173, out_174, out_175, out_176, out_177, out_178, out_179, out_180, out_181, out_182, out_183, out_184, out_185, out_186, out_187, out_188, out_189, out_190, out_191, out_192, out_193, out_194, out_195, out_196, out_197, out_198, out_199, out_200, out_201, out_202, out_203, out_204, out_205, out_206, out_207, out_208, out_209, out_210, out_211, out_212, out_213, out_214, out_215, out_216, out_217, out_218, out_219, out_220, out_221, out_222, out_223, out_224, out_225, out_226, out_227, out_228, out_229, out_230, out_231, out_232, out_233, out_234, out_235, out_236, out_237, out_238, out_239, out_240, out_241, out_242, out_243, out_244, out_245, out_246, out_247, out_248, out_249, out_250, out_251, out_252, out_253, out_254, out_255, out_256, out_257, out_258, out_259, out_260, out_261, out_262, out_263, out_264, out_265, out_266, out_267, out_268, out_269, out_270, out_271, out_272, out_273, out_274, out_275, out_276, out_277, out_278, out_279, out_280, out_281, out_282, out_283, out_284, out_285, out_286, out_287, out_288, out_289, out_290, out_291, out_292, out_293, out_294, out_295, out_296, out_297, out_298, out_299, out_300, out_301, out_302, out_303, out_304, out_305, out_306, out_307, out_308, out_309, out_310, out_311, out_312, out_313, out_314, out_315, out_316, out_317, out_318, out_319, out_320, out_321, out_322, out_323, out_324, out_325, out_326, out_327, out_328, out_329, out_330, out_331, out_332, out_333, out_334, out_335, out_336, out_337, out_338, out_339, out_340, out_341, out_342, out_343, out_344, out_345, out_346, out_347, out_348, out_349, out_350, out_351, out_352, out_353, out_354, out_355, out_356, out_357, out_358, out_359, out_360, out_361, out_362, out_363, out_364, out_365, out_366, out_367, out_368, out_369, out_370, out_371, out_372, out_373, out_374, out_375, out_376, out_377, out_378, out_379, out_380, out_381, out_382, out_383, out_384, out_385, out_386, out_387, out_388, out_389, out_390, out_391, out_392, out_393, out_394, out_395, out_396, out_397, out_398, out_399, out_400, out_401, out_402, out_403, out_404, out_405, out_406, out_407, out_408, out_409, out_410, out_411, out_412, out_413, out_414, out_415, out_416, out_417, out_418, out_419, out_420, out_421, out_422, out_423, out_424, out_425, out_426, out_427, out_428, out_429, out_430, out_431, out_432, out_433, out_434, out_435, out_436, out_437, out_438, out_439, out_440, out_441, out_442, out_443, out_444, out_445, out_446, out_447, out_448, out_449, out_450, out_451, out_452, out_453, out_454, out_455, out_456, out_457, out_458, out_459, out_460, out_461, out_462, out_463, out_464, out_465, out_466, out_467, out_468, out_469, out_470, out_471, out_472, out_473, out_474, out_475, out_476, out_477, out_478, out_479, out_480, out_481, out_482, out_483, out_484, out_485, out_486, out_487, out_488, out_489, out_490, out_491, out_492, out_493, out_494, out_495, out_496, out_497, out_498, out_499, out_500, out_501, out_502, out_503, out_504, out_505, out_506, out_507, out_508, out_509, out_510, out_511, out_512, out_513, out_514, out_515, out_516, out_517, out_518, out_519, out_520, out_521, out_522, out_523, out_524, out_525, out_526, out_527, out_528, out_529, out_530, out_531, out_532, out_533, out_534, out_535, out_536, out_537, out_538, out_539, out_540, out_541, out_542, out_543, out_544, out_545, out_546, out_547, out_548, out_549, out_550, out_551, out_552, out_553, out_554, out_555, out_556, out_557, out_558, out_559, out_560, out_561, out_562, out_563, out_564, out_565, out_566, out_567, out_568, out_569, out_570, out_571, out_572, out_573, out_574, out_575, out_576, out_577, out_578, out_579, out_580, out_581, out_582, out_583, out_584, out_585, out_586, out_587, out_588, out_589, out_590, out_591, out_592, out_593, out_594, out_595, out_596, out_597, out_598, out_599, out_600, out_601, out_602, out_603, out_604, out_605, out_606, out_607, out_608, out_609, out_610, out_611, out_612, out_613, out_614, out_615, out_616, out_617, out_618, out_619, out_620, out_621, out_622, out_623, out_624, out_625, out_626, out_627, out_628, out_629, out_630, out_631, out_632, out_633, out_634, out_635, out_636, out_637, out_638, out_639, out_640, out_641, out_642, out_643, out_644, out_645, out_646, out_647, out_648, out_649, out_650, out_651, out_652, out_653, out_654, out_655, out_656, out_657, out_658, out_659, out_660, out_661, out_662, out_663, out_664, out_665, out_666, out_667, out_668, out_669, out_670, out_671, out_672, out_673, out_674, out_675, out_676, out_677, out_678, out_679, out_680, out_681, out_682, out_683, out_684, out_685, out_686, out_687, out_688, out_689, out_690, out_691, out_692, out_693, out_694, out_695, out_696, out_697, out_698, out_699, out_700, out_701, out_702, out_703, out_704, out_705, out_706, out_707, out_708, out_709, out_710, out_711, out_712, out_713, out_714, out_715, out_716, out_717, out_718, out_719, out_720, out_721, out_722, out_723, out_724, out_725, out_726, out_727, out_728, out_729, out_730, out_731, out_732, out_733, out_734, out_735, out_736, out_737, out_738, out_739, out_740, out_741, out_742, out_743, out_744, out_745, out_746, out_747, out_748, out_749, out_750, out_751, out_752, out_753, out_754, out_755, out_756, out_757, out_758, out_759, out_760, out_761, out_762, out_763, out_764, out_765, out_766, out_767, out_768, out_769, out_770, out_771, out_772, out_773, out_774, out_775, out_776, out_777, out_778, out_779, out_780, out_781, out_782, out_783, out_784, out_785, out_786, out_787, out_788, out_789, out_790, out_791, out_792, out_793, out_794, out_795, out_796, out_797, out_798, out_799, out_800, out_801, out_802, out_803, out_804, out_805, out_806, out_807, out_808, out_809, out_810, out_811, out_812, out_813, out_814, out_815, out_816, out_817, out_818, out_819, out_820, out_821, out_822, out_823, out_824, out_825, out_826, out_827, out_828, out_829, out_830, out_831, out_832, out_833, out_834, out_835, out_836, out_837, out_838, out_839, out_840, out_841, out_842, out_843, out_844, out_845, out_846, out_847, out_848, out_849, out_850, out_851, out_852, out_853, out_854, out_855, out_856, out_857, out_858, out_859, out_860, out_861, out_862, out_863, out_864, out_865, out_866, out_867, out_868, out_869, out_870, out_871, out_872, out_873, out_874, out_875, out_876, out_877, out_878, out_879, out_880, out_881, out_882, out_883, out_884, out_885, out_886, out_887, out_888, out_889, out_890, out_891, out_892, out_893, out_894, out_895, out_896, out_897, out_898, out_899, out_900, out_901, out_902, out_903, out_904, out_905, out_906, out_907, out_908, out_909, out_910, out_911, out_912, out_913, out_914, out_915, out_916, out_917, out_918, out_919, out_920, out_921, out_922, out_923, out_924, out_925, out_926, out_927, out_928, out_929, out_930, out_931, out_932, out_933, out_934, out_935, out_936, out_937, out_938, out_939, out_940, out_941, out_942, out_943, out_944, out_945, out_946, out_947, out_948, out_949, out_950, out_951, out_952, out_953, out_954, out_955, out_956, out_957, out_958, out_959, out_960, out_961, out_962, out_963, out_964, out_965, out_966, out_967, out_968, out_969, out_970, out_971, out_972, out_973, out_974, out_975, out_976, out_977, out_978, out_979, out_980, out_981, out_982, out_983, out_984, out_985, out_986, out_987, out_988, out_989, out_990, out_991, out_992, out_993, out_994, out_995, out_996, out_997, out_998, out_999, out_1000, out_1001, out_1002, out_1003, out_1004, out_1005, out_1006, out_1007, out_1008, out_1009, out_1010, out_1011, out_1012, out_1013, out_1014, out_1015, out_1016, out_1017, out_1018, out_1019, out_1020, out_1021, out_1022, out_1023, out_1024, out_1025, out_1026, out_1027, out_1028, out_1029, out_1030, out_1031, out_1032, out_1033, out_1034, out_1035, out_1036, out_1037, out_1038, out_1039, out_1040, out_1041, out_1042, out_1043, out_1044, out_1045, out_1046, out_1047, out_1048, out_1049, out_1050, out_1051, out_1052, out_1053, out_1054, out_1055, out_1056, out_1057, out_1058, out_1059, out_1060, out_1061, out_1062, out_1063, out_1064, out_1065, out_1066, out_1067, out_1068, out_1069, out_1070, out_1071, out_1072, out_1073, out_1074, out_1075, out_1076, out_1077, out_1078, out_1079, out_1080, out_1081, out_1082, out_1083, out_1084, out_1085, out_1086, out_1087, out_1088, out_1089, out_1090, out_1091, out_1092, out_1093, out_1094, out_1095, out_1096, out_1097, out_1098, out_1099, out_1100, out_1101, out_1102, out_1103, out_1104, out_1105, out_1106, out_1107}, {out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[], out[0]});

fanout_n #(3, 0, 0) FANOUT_1 (maxAbsValueCir_wire_7, {maxAbsValueCir_wire_7_0, maxAbsValueCir_wire_7_1, maxAbsValueCir_wire_7_2});
fanout_n #(3, 0, 0) FANOUT_2 (maxAbsValueCir_wire_25, {maxAbsValueCir_wire_25_0, maxAbsValueCir_wire_25_1, maxAbsValueCir_wire_25_2});
fanout_n #(2, 0, 0) FANOUT_3 (maxAbsValueCir_wire_14, {maxAbsValueCir_wire_14_0, maxAbsValueCir_wire_14_1});
fanout_n #(2, 0, 0) FANOUT_4 (maxAbsValueCir_wire_5, {maxAbsValueCir_wire_5_0, maxAbsValueCir_wire_5_1});
fanout_n #(2, 0, 0) FANOUT_5 (maxAbsValueCir_wire_23, {maxAbsValueCir_wire_23_0, maxAbsValueCir_wire_23_1});
fanout_n #(8, 0, 0) FANOUT_6 (maxAbsValueCir_wire_57, {maxAbsValueCir_wire_57_0, maxAbsValueCir_wire_57_1, maxAbsValueCir_wire_57_2, maxAbsValueCir_wire_57_3, maxAbsValueCir_wire_57_4, maxAbsValueCir_wire_57_5, maxAbsValueCir_wire_57_6, maxAbsValueCir_wire_57_7});
fanout_n #(8, 0, 0) FANOUT_7 (maxAbsValueCir_wire_85, {maxAbsValueCir_wire_85_0, maxAbsValueCir_wire_85_1, maxAbsValueCir_wire_85_2, maxAbsValueCir_wire_85_3, maxAbsValueCir_wire_85_4, maxAbsValueCir_wire_85_5, maxAbsValueCir_wire_85_6, maxAbsValueCir_wire_85_7});
fanout_n #(4, 0, 0) FANOUT_8 (maxAbsValueCir_wire_59, {maxAbsValueCir_wire_59_0, maxAbsValueCir_wire_59_1, maxAbsValueCir_wire_59_2, maxAbsValueCir_wire_59_3});
fanout_n #(4, 0, 0) FANOUT_9 (maxAbsValueCir_wire_58, {maxAbsValueCir_wire_58_0, maxAbsValueCir_wire_58_1, maxAbsValueCir_wire_58_2, maxAbsValueCir_wire_58_3});
fanout_n #(6, 0, 0) FANOUT_10 (maxAbsValueCir_wire_34, {maxAbsValueCir_wire_34_0, maxAbsValueCir_wire_34_1, maxAbsValueCir_wire_34_2, maxAbsValueCir_wire_34_3, maxAbsValueCir_wire_34_4, maxAbsValueCir_wire_34_5});
fanout_n #(2, 0, 0) FANOUT_11 (maxAbsValueCir_wire_53, {maxAbsValueCir_wire_53_0, maxAbsValueCir_wire_53_1});
fanout_n #(2, 0, 0) FANOUT_12 (maxAbsValueCir_wire_44, {maxAbsValueCir_wire_44_0, maxAbsValueCir_wire_44_1});
fanout_n #(2, 0, 0) FANOUT_13 (maxAbsValueCir_wire_81, {maxAbsValueCir_wire_81_0, maxAbsValueCir_wire_81_1});
fanout_n #(2, 0, 0) FANOUT_14 (maxAbsValueCir_wire_72, {maxAbsValueCir_wire_72_0, maxAbsValueCir_wire_72_1});
fanout_n #(5, 0, 0) FANOUT_15 (maxAbsValueCir_wire_11, {maxAbsValueCir_wire_11_0, maxAbsValueCir_wire_11_1, maxAbsValueCir_wire_11_2, maxAbsValueCir_wire_11_3, maxAbsValueCir_wire_11_4});
fanout_n #(4, 0, 0) FANOUT_16 (maxAbsValueCir_wire_12, {maxAbsValueCir_wire_12_0, maxAbsValueCir_wire_12_1, maxAbsValueCir_wire_12_2, maxAbsValueCir_wire_12_3});
fanout_n #(4, 0, 0) FANOUT_17 (maxAbsValueCir_wire_15, {maxAbsValueCir_wire_15_0, maxAbsValueCir_wire_15_1, maxAbsValueCir_wire_15_2, maxAbsValueCir_wire_15_3});
fanout_n #(7, 0, 0) FANOUT_18 (maxAbsValueCir_wire_18, {maxAbsValueCir_wire_18_0, maxAbsValueCir_wire_18_1, maxAbsValueCir_wire_18_2, maxAbsValueCir_wire_18_3, maxAbsValueCir_wire_18_4, maxAbsValueCir_wire_18_5, maxAbsValueCir_wire_18_6});
fanout_n #(4, 0, 0) FANOUT_19 (maxAbsValueCir_wire_2, {maxAbsValueCir_wire_2_0, maxAbsValueCir_wire_2_1, maxAbsValueCir_wire_2_2, maxAbsValueCir_wire_2_3});
fanout_n #(4, 0, 0) FANOUT_20 (maxAbsValueCir_wire_3, {maxAbsValueCir_wire_3_0, maxAbsValueCir_wire_3_1, maxAbsValueCir_wire_3_2, maxAbsValueCir_wire_3_3});
fanout_n #(4, 0, 0) FANOUT_21 (maxAbsValueCir_wire_6, {maxAbsValueCir_wire_6_0, maxAbsValueCir_wire_6_1, maxAbsValueCir_wire_6_2, maxAbsValueCir_wire_6_3});
fanout_n #(9, 0, 0) FANOUT_22 (maxAbsValueCir_wire_9, {maxAbsValueCir_wire_9_0, maxAbsValueCir_wire_9_1, maxAbsValueCir_wire_9_2, maxAbsValueCir_wire_9_3, maxAbsValueCir_wire_9_4, maxAbsValueCir_wire_9_5, maxAbsValueCir_wire_9_6, maxAbsValueCir_wire_9_7, maxAbsValueCir_wire_9_8});
fanout_n #(4, 0, 0) FANOUT_23 (maxAbsValueCir_wire_20, {maxAbsValueCir_wire_20_0, maxAbsValueCir_wire_20_1, maxAbsValueCir_wire_20_2, maxAbsValueCir_wire_20_3});
fanout_n #(4, 0, 0) FANOUT_24 (maxAbsValueCir_wire_21, {maxAbsValueCir_wire_21_0, maxAbsValueCir_wire_21_1, maxAbsValueCir_wire_21_2, maxAbsValueCir_wire_21_3});
fanout_n #(4, 0, 0) FANOUT_25 (maxAbsValueCir_wire_24, {maxAbsValueCir_wire_24_0, maxAbsValueCir_wire_24_1, maxAbsValueCir_wire_24_2, maxAbsValueCir_wire_24_3});
fanout_n #(9, 0, 0) FANOUT_26 (maxAbsValueCir_wire_27, {maxAbsValueCir_wire_27_0, maxAbsValueCir_wire_27_1, maxAbsValueCir_wire_27_2, maxAbsValueCir_wire_27_3, maxAbsValueCir_wire_27_4, maxAbsValueCir_wire_27_5, maxAbsValueCir_wire_27_6, maxAbsValueCir_wire_27_7, maxAbsValueCir_wire_27_8});


xor_n #(2, 0, 0) XOR_1 (maxAbsValueCir_wire_1, {maxAbsValueCir_wire_2_0, maxAbsValueCir_wire_3_0});
xnor_n #(2, 0, 0) XNOR_1 (maxAbsValueCir_wire_4, {maxAbsValueCir_wire_5_0, maxAbsValueCir_wire_6_0});
xnor_n #(2, 0, 0) XNOR_2 (maxAbsValueCir_wire_7, {maxAbsValueCir_wire_8, maxAbsValueCir_wire_9_0});
xor_n #(2, 0, 0) XOR_2 (maxAbsValueCir_wire_10, {maxAbsValueCir_wire_11_0, maxAbsValueCir_wire_12_0});
xnor_n #(2, 0, 0) XNOR_3 (maxAbsValueCir_wire_13, {maxAbsValueCir_wire_14_0, maxAbsValueCir_wire_15_0});
xnor_n #(2, 0, 0) XNOR_4 (maxAbsValueCir_wire_16, {maxAbsValueCir_wire_17, maxAbsValueCir_wire_18_0});
xor_n #(2, 0, 0) XOR_3 (maxAbsValueCir_wire_19, {maxAbsValueCir_wire_20_0, maxAbsValueCir_wire_21_0});
xnor_n #(2, 0, 0) XNOR_5 (maxAbsValueCir_wire_22, {maxAbsValueCir_wire_23_0, maxAbsValueCir_wire_24_0});
xnor_n #(2, 0, 0) XNOR_6 (maxAbsValueCir_wire_25, {maxAbsValueCir_wire_26, maxAbsValueCir_wire_27_0});
and_n #(2, 0, 0) AND_1 (maxAbsValueCir_wire_17, {maxAbsValueCir_wire_14_1, maxAbsValueCir_wire_28});
nor_n #(2, 0, 0) NOR_1 (maxAbsValueCir_wire_14, {maxAbsValueCir_wire_12_1, maxAbsValueCir_wire_11_1});
notg #(0, 0) NOT_1 (maxAbsValueCir_wire_28, maxAbsValueCir_wire_15_1);
and_n #(2, 0, 0) AND_2 (maxAbsValueCir_wire_8, {maxAbsValueCir_wire_5_1, maxAbsValueCir_wire_29});
nor_n #(2, 0, 0) NOR_2 (maxAbsValueCir_wire_5, {maxAbsValueCir_wire_3_1, maxAbsValueCir_wire_2_1});
notg #(0, 0) NOT_2 (maxAbsValueCir_wire_29, maxAbsValueCir_wire_6_1);
and_n #(2, 0, 0) AND_3 (maxAbsValueCir_wire_26, {maxAbsValueCir_wire_23_1, maxAbsValueCir_wire_30});
nor_n #(2, 0, 0) NOR_3 (maxAbsValueCir_wire_23, {maxAbsValueCir_wire_21_1, maxAbsValueCir_wire_20_1});
notg #(0, 0) NOT_3 (maxAbsValueCir_wire_30, maxAbsValueCir_wire_24_1);
and_n #(2, 0, 0) AND_4 (maxAbsValueCir_wire_31, {maxAbsValueCir_wire_7_0, maxAbsValueCir_wire_9_1});
and_n #(2, 0, 0) AND_5 (maxAbsValueCir_wire_32, {maxAbsValueCir_wire_31, maxAbsValueCir_wire_33});
notg #(0, 0) NOT_4 (maxAbsValueCir_wire_33, maxAbsValueCir_wire_34_0);
notg #(0, 0) NOT_5 (maxAbsValueCir_wire_35, maxAbsValueCir_wire_11_2);
and_n #(3, 0, 0) AND_6 (maxAbsValueCir_wire_36, {maxAbsValueCir_wire_35, maxAbsValueCir_wire_37, maxAbsValueCir_wire_2_2});
or_n #(2, 0, 0) OR_1 (maxAbsValueCir_wire_38, {maxAbsValueCir_wire_32, maxAbsValueCir_wire_39});
or_n #(2, 0, 0) OR_2 (maxAbsValueCir_wire_40, {maxAbsValueCir_wire_41, maxAbsValueCir_wire_42});
and_n #(3, 0, 0) AND_7 (maxAbsValueCir_wire_39, {maxAbsValueCir_wire_40, maxAbsValueCir_wire_43, maxAbsValueCir_wire_44_0});
or_n #(2, 0, 0) OR_3 (maxAbsValueCir_wire_45, {maxAbsValueCir_wire_46, maxAbsValueCir_wire_44_1});
and_n #(2, 0, 0) AND_8 (maxAbsValueCir_wire_47, {maxAbsValueCir_wire_45, maxAbsValueCir_wire_48});
or_n #(2, 0, 0) OR_4 (maxAbsValueCir_wire_48, {maxAbsValueCir_wire_49, maxAbsValueCir_wire_50});
and_n #(2, 0, 0) AND_9 (maxAbsValueCir_wire_51, {maxAbsValueCir_wire_52, maxAbsValueCir_wire_53_0});
or_n #(2, 0, 0) OR_5 (maxAbsValueCir_wire_54, {maxAbsValueCir_wire_51, maxAbsValueCir_wire_36});
or_n #(2, 0, 0) OR_6 (maxAbsValueCir_wire_37, {maxAbsValueCir_wire_55, maxAbsValueCir_wire_53_1});
and_n #(2, 0, 0) AND_10 (maxAbsValueCir_wire_56, {maxAbsValueCir_wire_47, maxAbsValueCir_wire_54});
and_n #(2, 0, 0) AND_11 (maxAbsValueCir_wire_41, {maxAbsValueCir_wire_7_1, maxAbsValueCir_wire_9_2});
or_n #(2, 0, 0) OR_7 (maxAbsValueCir_wire_57, {maxAbsValueCir_wire_38, maxAbsValueCir_wire_56});
notg #(0, 0) NOT_6 (maxAbsValueCir_wire_42, maxAbsValueCir_wire_34_1);
notg #(0, 0) NOT_7 (maxAbsValueCir_wire_43, maxAbsValueCir_wire_58_0);
notg #(0, 0) NOT_8 (maxAbsValueCir_wire_46, maxAbsValueCir_wire_58_1);
and_n #(2, 0, 0) AND_12 (maxAbsValueCir_wire_49, {maxAbsValueCir_wire_7_2, maxAbsValueCir_wire_9_3});
notg #(0, 0) NOT_9 (maxAbsValueCir_wire_50, maxAbsValueCir_wire_34_2);
notg #(0, 0) NOT_10 (maxAbsValueCir_wire_52, maxAbsValueCir_wire_59_0);
notg #(0, 0) NOT_11 (maxAbsValueCir_wire_55, maxAbsValueCir_wire_59_1);
and_n #(2, 0, 0) AND_13 (maxAbsValueCir_wire_60, {maxAbsValueCir_wire_25_0, maxAbsValueCir_wire_27_1});
and_n #(2, 0, 0) AND_14 (maxAbsValueCir_wire_61, {maxAbsValueCir_wire_60, maxAbsValueCir_wire_62});
notg #(0, 0) NOT_12 (maxAbsValueCir_wire_62, maxAbsValueCir_wire_34_3);
notg #(0, 0) NOT_13 (maxAbsValueCir_wire_63, maxAbsValueCir_wire_11_3);
and_n #(3, 0, 0) AND_15 (maxAbsValueCir_wire_64, {maxAbsValueCir_wire_63, maxAbsValueCir_wire_65, maxAbsValueCir_wire_20_2});
or_n #(2, 0, 0) OR_8 (maxAbsValueCir_wire_66, {maxAbsValueCir_wire_61, maxAbsValueCir_wire_67});
or_n #(2, 0, 0) OR_9 (maxAbsValueCir_wire_68, {maxAbsValueCir_wire_69, maxAbsValueCir_wire_70});
and_n #(3, 0, 0) AND_16 (maxAbsValueCir_wire_67, {maxAbsValueCir_wire_68, maxAbsValueCir_wire_71, maxAbsValueCir_wire_72_0});
or_n #(2, 0, 0) OR_10 (maxAbsValueCir_wire_73, {maxAbsValueCir_wire_74, maxAbsValueCir_wire_72_1});
and_n #(2, 0, 0) AND_17 (maxAbsValueCir_wire_75, {maxAbsValueCir_wire_73, maxAbsValueCir_wire_76});
or_n #(2, 0, 0) OR_11 (maxAbsValueCir_wire_76, {maxAbsValueCir_wire_77, maxAbsValueCir_wire_78});
and_n #(2, 0, 0) AND_18 (maxAbsValueCir_wire_79, {maxAbsValueCir_wire_80, maxAbsValueCir_wire_81_0});
or_n #(2, 0, 0) OR_12 (maxAbsValueCir_wire_82, {maxAbsValueCir_wire_79, maxAbsValueCir_wire_64});
or_n #(2, 0, 0) OR_13 (maxAbsValueCir_wire_65, {maxAbsValueCir_wire_83, maxAbsValueCir_wire_81_1});
and_n #(2, 0, 0) AND_19 (maxAbsValueCir_wire_84, {maxAbsValueCir_wire_75, maxAbsValueCir_wire_82});
and_n #(2, 0, 0) AND_20 (maxAbsValueCir_wire_69, {maxAbsValueCir_wire_25_1, maxAbsValueCir_wire_27_2});
or_n #(2, 0, 0) OR_14 (maxAbsValueCir_wire_85, {maxAbsValueCir_wire_66, maxAbsValueCir_wire_84});
notg #(0, 0) NOT_14 (maxAbsValueCir_wire_70, maxAbsValueCir_wire_34_4);
notg #(0, 0) NOT_15 (maxAbsValueCir_wire_71, maxAbsValueCir_wire_58_2);
notg #(0, 0) NOT_16 (maxAbsValueCir_wire_74, maxAbsValueCir_wire_58_3);
and_n #(2, 0, 0) AND_21 (maxAbsValueCir_wire_77, {maxAbsValueCir_wire_25_2, maxAbsValueCir_wire_27_3});
notg #(0, 0) NOT_17 (maxAbsValueCir_wire_78, maxAbsValueCir_wire_34_5);
notg #(0, 0) NOT_18 (maxAbsValueCir_wire_80, maxAbsValueCir_wire_59_2);
notg #(0, 0) NOT_19 (maxAbsValueCir_wire_83, maxAbsValueCir_wire_59_3);
or_n #(2, 0, 0) OR_15 (maxAbsValueCir_wire_59, {maxAbsValueCir_wire_86, maxAbsValueCir_wire_87});
and_n #(2, 0, 0) AND_22 (maxAbsValueCir_wire_86, {maxAbsValueCir_wire_10, maxAbsValueCir_wire_18_1});
notg #(0, 0) NOT_20 (maxAbsValueCir_wire_88, maxAbsValueCir_wire_18_2);
and_n #(2, 0, 0) AND_23 (maxAbsValueCir_wire_87, {maxAbsValueCir_wire_88, maxAbsValueCir_wire_12_2});
or_n #(2, 0, 0) OR_16 (maxAbsValueCir_wire_58, {maxAbsValueCir_wire_89, maxAbsValueCir_wire_90});
and_n #(2, 0, 0) AND_24 (maxAbsValueCir_wire_89, {maxAbsValueCir_wire_13, maxAbsValueCir_wire_18_3});
notg #(0, 0) NOT_21 (maxAbsValueCir_wire_91, maxAbsValueCir_wire_18_4);
and_n #(2, 0, 0) AND_25 (maxAbsValueCir_wire_90, {maxAbsValueCir_wire_91, maxAbsValueCir_wire_15_2});
and_n #(2, 0, 0) AND_26 (maxAbsValueCir_wire_34, {maxAbsValueCir_wire_16, maxAbsValueCir_wire_18_5});
or_n #(2, 0, 0) OR_17 (maxAbsValueCir_wire_53, {maxAbsValueCir_wire_92, maxAbsValueCir_wire_93});
and_n #(2, 0, 0) AND_27 (maxAbsValueCir_wire_92, {maxAbsValueCir_wire_1, maxAbsValueCir_wire_9_4});
notg #(0, 0) NOT_22 (maxAbsValueCir_wire_94, maxAbsValueCir_wire_9_5);
and_n #(2, 0, 0) AND_28 (maxAbsValueCir_wire_93, {maxAbsValueCir_wire_94, maxAbsValueCir_wire_3_2});
or_n #(2, 0, 0) OR_18 (maxAbsValueCir_wire_44, {maxAbsValueCir_wire_95, maxAbsValueCir_wire_96});
and_n #(2, 0, 0) AND_29 (maxAbsValueCir_wire_95, {maxAbsValueCir_wire_4, maxAbsValueCir_wire_9_6});
notg #(0, 0) NOT_23 (maxAbsValueCir_wire_97, maxAbsValueCir_wire_9_7);
and_n #(2, 0, 0) AND_30 (maxAbsValueCir_wire_96, {maxAbsValueCir_wire_97, maxAbsValueCir_wire_6_2});
or_n #(2, 0, 0) OR_19 (maxAbsValueCir_wire_81, {maxAbsValueCir_wire_98, maxAbsValueCir_wire_99});
and_n #(2, 0, 0) AND_31 (maxAbsValueCir_wire_98, {maxAbsValueCir_wire_19, maxAbsValueCir_wire_27_4});
notg #(0, 0) NOT_24 (maxAbsValueCir_wire_100, maxAbsValueCir_wire_27_5);
and_n #(2, 0, 0) AND_32 (maxAbsValueCir_wire_99, {maxAbsValueCir_wire_100, maxAbsValueCir_wire_21_2});
or_n #(2, 0, 0) OR_20 (maxAbsValueCir_wire_72, {maxAbsValueCir_wire_101, maxAbsValueCir_wire_102});
and_n #(2, 0, 0) AND_33 (maxAbsValueCir_wire_101, {maxAbsValueCir_wire_22, maxAbsValueCir_wire_27_6});
notg #(0, 0) NOT_25 (maxAbsValueCir_wire_103, maxAbsValueCir_wire_27_7);
and_n #(2, 0, 0) AND_34 (maxAbsValueCir_wire_102, {maxAbsValueCir_wire_103, maxAbsValueCir_wire_24_2});
bufg #(0, 0) BUF_1 (out_3, maxAbsValueCir_wire_104);
and_n #(2, 0, 0) AND_35 (maxAbsValueCir_wire_105, {maxAbsValueCir_wire_57_0, maxAbsValueCir_wire_2_3});
or_n #(2, 0, 0) OR_21 (maxAbsValueCir_wire_104, {maxAbsValueCir_wire_105, maxAbsValueCir_wire_106});
and_n #(2, 0, 0) AND_36 (maxAbsValueCir_wire_107, {maxAbsValueCir_wire_85_0, maxAbsValueCir_wire_20_3});
or_n #(2, 0, 0) OR_22 (maxAbsValueCir_wire_108, {maxAbsValueCir_wire_107, maxAbsValueCir_wire_109});
notg #(0, 0) NOT_26 (maxAbsValueCir_wire_110, maxAbsValueCir_wire_85_1);
and_n #(2, 0, 0) AND_37 (maxAbsValueCir_wire_109, {maxAbsValueCir_wire_110, maxAbsValueCir_wire_11_4});
notg #(0, 0) NOT_27 (maxAbsValueCir_wire_111, maxAbsValueCir_wire_57_1);
and_n #(2, 0, 0) AND_38 (maxAbsValueCir_wire_106, {maxAbsValueCir_wire_111, maxAbsValueCir_wire_108});
bufg #(0, 0) BUF_2 (out_2, maxAbsValueCir_wire_112);
and_n #(2, 0, 0) AND_39 (maxAbsValueCir_wire_113, {maxAbsValueCir_wire_57_2, maxAbsValueCir_wire_3_3});
or_n #(2, 0, 0) OR_23 (maxAbsValueCir_wire_112, {maxAbsValueCir_wire_113, maxAbsValueCir_wire_114});
and_n #(2, 0, 0) AND_40 (maxAbsValueCir_wire_115, {maxAbsValueCir_wire_85_2, maxAbsValueCir_wire_21_3});
or_n #(2, 0, 0) OR_24 (maxAbsValueCir_wire_116, {maxAbsValueCir_wire_115, maxAbsValueCir_wire_117});
notg #(0, 0) NOT_28 (maxAbsValueCir_wire_118, maxAbsValueCir_wire_85_3);
and_n #(2, 0, 0) AND_41 (maxAbsValueCir_wire_117, {maxAbsValueCir_wire_118, maxAbsValueCir_wire_12_3});
notg #(0, 0) NOT_29 (maxAbsValueCir_wire_119, maxAbsValueCir_wire_57_3);
and_n #(2, 0, 0) AND_42 (maxAbsValueCir_wire_114, {maxAbsValueCir_wire_119, maxAbsValueCir_wire_116});
bufg #(0, 0) BUF_3 (out_1, maxAbsValueCir_wire_120);
and_n #(2, 0, 0) AND_43 (maxAbsValueCir_wire_121, {maxAbsValueCir_wire_57_4, maxAbsValueCir_wire_6_3});
or_n #(2, 0, 0) OR_25 (maxAbsValueCir_wire_120, {maxAbsValueCir_wire_121, maxAbsValueCir_wire_122});
and_n #(2, 0, 0) AND_44 (maxAbsValueCir_wire_123, {maxAbsValueCir_wire_85_4, maxAbsValueCir_wire_24_3});
or_n #(2, 0, 0) OR_26 (maxAbsValueCir_wire_124, {maxAbsValueCir_wire_123, maxAbsValueCir_wire_125});
notg #(0, 0) NOT_30 (maxAbsValueCir_wire_126, maxAbsValueCir_wire_85_5);
and_n #(2, 0, 0) AND_45 (maxAbsValueCir_wire_125, {maxAbsValueCir_wire_126, maxAbsValueCir_wire_15_3});
notg #(0, 0) NOT_31 (maxAbsValueCir_wire_127, maxAbsValueCir_wire_57_5);
and_n #(2, 0, 0) AND_46 (maxAbsValueCir_wire_122, {maxAbsValueCir_wire_127, maxAbsValueCir_wire_124});
bufg #(0, 0) BUF_4 (out_0, maxAbsValueCir_wire_128);
and_n #(2, 0, 0) AND_47 (maxAbsValueCir_wire_129, {maxAbsValueCir_wire_57_6, maxAbsValueCir_wire_9_8});
or_n #(2, 0, 0) OR_27 (maxAbsValueCir_wire_128, {maxAbsValueCir_wire_129, maxAbsValueCir_wire_130});
and_n #(2, 0, 0) AND_48 (maxAbsValueCir_wire_131, {maxAbsValueCir_wire_85_6, maxAbsValueCir_wire_27_8});
or_n #(2, 0, 0) OR_28 (maxAbsValueCir_wire_132, {maxAbsValueCir_wire_131, maxAbsValueCir_wire_133});
notg #(0, 0) NOT_32 (maxAbsValueCir_wire_134, maxAbsValueCir_wire_85_7);
and_n #(2, 0, 0) AND_49 (maxAbsValueCir_wire_133, {maxAbsValueCir_wire_134, maxAbsValueCir_wire_18_6});
notg #(0, 0) NOT_33 (maxAbsValueCir_wire_135, maxAbsValueCir_wire_57_7);
and_n #(2, 0, 0) AND_50 (maxAbsValueCir_wire_130, {maxAbsValueCir_wire_135, maxAbsValueCir_wire_132});
bufg #(0, 0) BUF_5 (maxAbsValueCir_wire_11, w1_3);
bufg #(0, 0) BUF_6 (maxAbsValueCir_wire_12, w1_2);
bufg #(0, 0) BUF_7 (maxAbsValueCir_wire_15, w1_1);
bufg #(0, 0) BUF_8 (maxAbsValueCir_wire_18, w1_0);
bufg #(0, 0) BUF_9 (maxAbsValueCir_wire_2, w2_3);
bufg #(0, 0) BUF_10 (maxAbsValueCir_wire_3, w2_2);
bufg #(0, 0) BUF_11 (maxAbsValueCir_wire_6, w2_1);
bufg #(0, 0) BUF_12 (maxAbsValueCir_wire_9, w2_0);
bufg #(0, 0) BUF_13 (maxAbsValueCir_wire_20, w3_3);
bufg #(0, 0) BUF_14 (maxAbsValueCir_wire_21, w3_2);
bufg #(0, 0) BUF_15 (maxAbsValueCir_wire_24, w3_1);
bufg #(0, 0) BUF_16 (maxAbsValueCir_wire_27, w3_0);

endmodule
