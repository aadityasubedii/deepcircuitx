    always @(posedge clk) begin
        divider <= divider + 1;
    end