always @(next_state) begin
	state = next_state; 
end