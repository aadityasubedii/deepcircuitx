    always @(negedge dqs_in[ 7]) dqs_neg_timing_check( 7);