always @ ( posedge reset, posedge clk ) begin
	if (reset) begin
		o_copro_read_data <= 'd0;
	end else begin       
	    if ( !i_core_stall )
		  case ( i_copro_crn )
		      
		      4'd0:    o_copro_read_data <= 32'h4156_0300;
		      4'd2:    o_copro_read_data <= {29'd0, cache_control}; 
		      4'd3:    o_copro_read_data <= cacheable_area; 
		      4'd4:    o_copro_read_data <= updateable_area; 
		      4'd5:    o_copro_read_data <= disruptive_area; 
		      4'd6:    o_copro_read_data <= {24'd0, fault_status };
		      4'd7:    o_copro_read_data <= fault_address;
		      default: o_copro_read_data <= 32'd0;
		  endcase
	end
end