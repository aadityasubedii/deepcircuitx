module KURM_controller(Out0, Out1, Out2, Out3, Out4, Out5A, Out5B, Out5C, Out5Active, Out6, Out7, Out8, s0, s1, s2, s3, clock);   

input s0, s1, s2, s3;
input clock;
output Out0,  Out1,  Out2,  Out3, Out4,  Out5A, Out5B, Out5C, Out5Active, Out6, Out7, Out8;















reg  out0,  out1,  out2,  out3, out4, out5A, out5B, out5C, out5Active, out6,  out7, out8;