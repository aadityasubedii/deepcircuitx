    always @(negedge dqs_in[11]) dqs_neg_timing_check(11);