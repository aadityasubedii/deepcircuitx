always @(posedge clk)
	b <= a;
