always @(posedge clock)    
begin
	
	tempA=registers[instructionAdd];
	
end