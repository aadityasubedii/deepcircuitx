  always @* begin
    
    $display("CLOCKS_PER_TICK: %d", CLOCKS_PER_TICK);
    $display("TICK_WIDTH: %d", TICK_WIDTH);
  end