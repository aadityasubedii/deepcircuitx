always@(posedge clk)
begin
	
		IN[0] <= DATA_IN;
		IN[1] <= IN[0];
		IN[2] <= IN[1];
		IN[3] <= IN[2];
		IN[4] <= IN[3];
		IN[5] <= IN[4];
		IN[6] <= IN[5];
		IN[7] <= IN[6];
		IN[8] <= IN[7];
		IN[9] <= IN[8];
		IN[10] <= IN[9];
		IN[11] <= IN[10];
		IN[12] <= IN[11];
		IN[13] <= IN[12];
		IN[14] <= IN[13];
		IN[15] <= IN[14];
		IN[16] <= IN[15];
		IN[17] <= IN[16];
		IN[18] <= IN[17];
		IN[19] <= IN[18];
		IN[20] <= IN[19];
		IN[21] <= IN[20];
        IN[22] <= IN[21];
        IN[23] <= IN[22];
        IN[24] <= IN[23];
        IN[25] <= IN[24];
        IN[26] <= IN[25];
        IN[27] <= IN[26];
        IN[28] <= IN[27];
        IN[29] <= IN[28];
        IN[30] <= IN[29];
        IN[31] <= IN[30];
        IN[32] <= IN[31];
        IN[33] <= IN[32];
        IN[34] <= IN[33];
        IN[35] <= IN[34];
        IN[36] <= IN[35];
        IN[37] <= IN[36];
        IN[38] <= IN[37];
        IN[39] <= IN[38];
        IN[40] <= IN[39];

end