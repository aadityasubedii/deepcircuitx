    always @(ck_n   ) ck_n_in    <= #BUS_DELAY ck_n;