    always @(posedge clk) sync_access <= !ce_n;