    always @(addr[3]) addr_timing_check(3);