    always @(dq_in[61]) dq_timing_check(61);