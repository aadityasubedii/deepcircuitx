            always @(posedge pll_ck) begin
                scale <= scale + 1;
            end