   always @(posedge clk)
			state <= nextstate;

   