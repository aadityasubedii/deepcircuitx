    always @(posedge dqs_even[ 8]) dqs_even_receiver( 8);