always @(posedge CLOCK_50) xck++;
