        always @* begin
            out_valid   = internal_out_valid;
            out_payload = internal_out_payload;
        end