always@ (UBn, Bn) begin
	
	BnP <= Bn + UBn;
end