        always @* begin
            fill_level = 0;
        end  