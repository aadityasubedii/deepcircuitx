    always @(posedge ck) begin
        out <= a * b;
    end