    always @(dq_in[46]) dq_timing_check(46);