  always @(posedge clk or negedge reset_n)