always @(A1,A1S) begin
	if (!A1S)
		FA1 <= (A1<=8191)?{A1[14:0], 2'b00}:(32764);
	else
		FA1 <= (A1>=57345)? {A1[14:0], 2'b00}: (98308);
end