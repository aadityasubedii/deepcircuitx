    always @(posedge ck) begin
        negative <= neg_audio;
    end