    always @(posedge ck) begin
        sck0 <= sck;
        ws0  <= ws;
    end