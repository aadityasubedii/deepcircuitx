always @(posedge clk)
	cur_test_clk	<= test_clk;
