always @(posedge clk)
	last_test_clk	<= cur_test_clk;
