module lab7_soc_nios2_gen2_0_cpu_nios2_oci_td_mode (
                                                     
                                                      ctrl,

                                                     
                                                      td_mode
                                                   )
;