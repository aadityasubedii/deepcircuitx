    always @(posedge ck) begin
        gain_0 <= gain;
    end