    always @(posedge mclk)begin
        r_cnt256_n <= r_cnt256_n - 8'd1;
    end