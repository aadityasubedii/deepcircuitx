    always @(ba_in  [ 0]) cmd_addr_timing_check( 4);