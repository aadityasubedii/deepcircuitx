module filter3(input clock,
                input signed [W-1:0]Xin,
                output reg signed [W-1:0]Y);