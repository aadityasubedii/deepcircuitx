module lab7_soc_jtag_uart_0_sim_scfifo_r (
                                           
                                            clk,
                                            fifo_rd,
                                            rst_n,

                                           
                                            fifo_EF,
                                            fifo_rdata,
                                            rfifo_full,
                                            rfifo_used
                                         )
;