    always @(posedge ck) begin
        prev_ws <= ws0;
        prev_sck <= sck0;
    end    