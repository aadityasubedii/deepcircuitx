always@ (MAG) begin

	casez (MAG)	
		15'b1??????????????:
			begin
				EXP <= 15;
			end
		15'b01?????????????:
			begin
				EXP <= 14;
			end
		15'b001????????????:
			begin
				EXP <= 13;
			end
		15'b0001???????????:
			begin
				EXP <= 12;
			end
		15'b00001??????????:
			begin
				EXP <= 11;
			end
		15'b000001?????????:
			begin
				EXP <= 10;
			end
		15'b0000001????????:
			begin
				EXP <= 9;
			end
		15'b00000001???????:
			begin
				EXP <= 8;
			end
		15'b000000001??????:
			begin
				EXP <= 7;
			end
		15'b0000000001?????:
			begin
				EXP <= 6;
			end
		15'b00000000001????:
			begin
				EXP <= 5;
			end
		15'b000000000001???:
			begin
				EXP <= 4;
			end
		15'b0000000000001??:
			begin
				EXP <= 3;
			end
		15'b00000000000001?:
			begin
				EXP <= 2;
			end
		15'b000000000000001:
			begin
				EXP <= 1;
			end
		default:
			begin
				EXP <= 0;
			end
	endcase
end