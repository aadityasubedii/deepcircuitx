        initial
            $display("Boot mem file is %s", `BOOT_MEM32_PARAMS_FILE );
    `endif
`endif

    
endmodule