always @(In1,In2)
begin
	temp=$signed(In1)+$signed(In2);
end