    always @(dq_in[39]) dq_timing_check(39);