			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end