    always @(posedge dqs_in[ 8]) dqs_pos_timing_check( 8);