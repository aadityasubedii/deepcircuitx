            always @(posedge ck) begin
                reseter <= reseter + 1;
            end