always @(posedge AUD_BCLK) sync <= AUD_DACLRCK;