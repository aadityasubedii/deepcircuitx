module pll(
    input wire clock_in,
    output wire clock_out,
    output wire locked
);