        always @* begin
            reset_out = reset_out_pre2;
            reset_req = reset_req_pre;
        end