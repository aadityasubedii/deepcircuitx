    always @(addr[2]) addr_timing_check(2);