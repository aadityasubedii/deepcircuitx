module fsm_reaction(
	clk,
	tick,
	trigger,
	time_out,
	count_over,
	en_lfsr,
	start_delay,
	start_count,
	reset_count,
	ledr
);