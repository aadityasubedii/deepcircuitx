assign dataOut=tempA;    
	
endmodule