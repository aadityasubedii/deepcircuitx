module C_LUT // #(.data_size(xx)) 
(
  input   [11:0]  step_counter,
  output  [15:0]  wave
);
always @(step_counter)
begin
  case(step_counter)
    1   : wave = 32624;
    2   : wave = 32380;
    3   : wave = 32542;
    4   : wave = 32629;
    5   : wave = 32479;
    6   : wave = 32325;
    7   : wave = 32484;
    8   : wave = 32731;
    9   : wave = 32661;
    10  : wave = 32815;
    11  : wave = 32621;
    12  : wave = 32588;
    13  : wave = 32670;
    14  : wave = 32655;
    15  : wave = 32830;
    16  : wave = 32827;
    17  : wave = 32771;
    18  : wave = 32835;
    19  : wave = 32876;
    20  : wave = 32958;
    21  : wave = 33088;
    22  : wave = 33042;
    23  : wave = 33084;
    24  : wave = 33029;
    25  : wave = 33050;
    26  : wave = 32809;
    27  : wave = 32768;
    28  : wave = 33044;
    29  : wave = 33068;
    30  : wave = 32977;
    31  : wave = 32919;
    32  : wave = 33062;
    33  : wave = 33206;
    34  : wave = 33160;
    35  : wave = 33258;
    36  : wave = 33830;
    37  : wave = 33448;
    38  : wave = 34098;
    39  : wave = 33657;
    40  : wave = 37675;
    41  : wave = 47525;
    42  : wave = 44215;
    43  : wave = 35444;
    44  : wave = 35762;
    45  : wave = 38607;
    46  : wave = 41007;
    47  : wave = 41464;
    48  : wave = 37823;
    49  : wave = 35430;
    50  : wave = 35098;
    51  : wave = 35859;
    52  : wave = 40693;
    53  : wave = 42268;
    54  : wave = 36598;
    55  : wave = 26454;
    56  : wave = 21206;
    57  : wave = 24894;
    58  : wave = 27302;
    59  : wave = 25245;
    60  : wave = 22047;
    61  : wave = 20726;
    62  : wave = 19812;
    63  : wave = 20744;
    64  : wave = 24961;
    65  : wave = 26071;
    66  : wave = 19302;
    67  : wave = 11837;
    68  : wave = 13902;
    69  : wave = 21327;
    70  : wave = 26554;
    71  : wave = 26983;
    72  : wave = 25549;
    73  : wave = 26910;
    74  : wave = 29716;
    75  : wave = 31245;
    76  : wave = 32179;
    77  : wave = 33499;
    78  : wave = 31681;
    79  : wave = 29519;
    80  : wave = 32873;
    81  : wave = 37329;
    82  : wave = 40309;
    83  : wave = 41041;
    84  : wave = 39311;
    85  : wave = 38137;
    86  : wave = 36578;
    87  : wave = 35557;
    88  : wave = 35852;
    89  : wave = 35066;
    90  : wave = 32676;
    91  : wave = 31126;
    92  : wave = 32008;
    93  : wave = 33271;
    94  : wave = 33041;
    95  : wave = 30827;
    96  : wave = 30973;
    97  : wave = 35096;
    98  : wave = 34983;
    99  : wave = 34156;
    100 : wave = 37518;
    101 : wave = 33375;
    102 : wave = 30230;
    103 : wave = 37011;
    104 : wave = 36405;
    105 : wave = 33963;
    106 : wave = 38081;
    107 : wave = 37419;
    108 : wave = 38673;
    109 : wave = 42817;
    110 : wave = 40129;
    111 : wave = 37367;
    112 : wave = 37348;
    113 : wave = 35139;
    114 : wave = 31584;
    115 : wave = 30117;
    116 : wave = 31126;
    117 : wave = 31906;
    118 : wave = 31021;
    119 : wave = 30436;
    120 : wave = 30705;
    121 : wave = 30906;
    122 : wave = 28686;
    123 : wave = 26869;
    124 : wave = 26396;
    125 : wave = 21955;
    126 : wave = 24456;
    127 : wave = 29554;
    128 : wave = 28900;
    129 : wave = 32757;
    130 : wave = 33279;
    131 : wave = 30592;
    132 : wave = 33662;
    133 : wave = 33737;
    134 : wave = 30781;
    135 : wave = 32864;
    136 : wave = 33178;
    137 : wave = 32417;
    138 : wave = 36683;
    139 : wave = 38154;
    140 : wave = 38322;
    141 : wave = 40528;
    142 : wave = 37652;
    143 : wave = 33651;
    144 : wave = 33959;
    145 : wave = 32241;
    146 : wave = 31900;
    147 : wave = 34683;
    148 : wave = 32348;
    149 : wave = 31007;
    150 : wave = 34689;
    151 : wave = 34489;
    152 : wave = 32359;
    153 : wave = 30889;
    154 : wave = 26130;
    155 : wave = 26315;
    156 : wave = 30419;
    157 : wave = 28297;
    158 : wave = 28996;
    159 : wave = 32183;
    160 : wave = 32214;
    161 : wave = 34075;
    162 : wave = 30703;
    163 : wave = 28507;
    164 : wave = 33496;
    165 : wave = 33592;
    166 : wave = 30734;
    167 : wave = 32701;
    168 : wave = 37300;
    169 : wave = 38398;
    170 : wave = 38557;
    171 : wave = 37806;
    172 : wave = 37287;
    173 : wave = 37736;
    174 : wave = 34909;
    175 : wave = 34501;
    176 : wave = 36903;
    177 : wave = 36555;
    178 : wave = 35525;
    179 : wave = 39100;
    180 : wave = 40318;
    181 : wave = 37756;
    182 : wave = 36767;
    183 : wave = 33747;
    184 : wave = 32597;
    185 : wave = 31785;
    186 : wave = 31526;
    187 : wave = 34373;
    188 : wave = 34327;
    189 : wave = 36756;
    190 : wave = 37977;
    191 : wave = 33480;
    192 : wave = 35899;
    193 : wave = 36676;
    194 : wave = 29943;
    195 : wave = 31483;
    196 : wave = 32627;
    197 : wave = 29711;
    198 : wave = 34716;
    199 : wave = 37434;
    200 : wave = 36096;
    201 : wave = 36987;
    202 : wave = 36566;
    203 : wave = 33851;
    204 : wave = 33580;
    205 : wave = 35121;
    206 : wave = 31799;
    207 : wave = 33312;
    208 : wave = 35777;
    209 : wave = 33016;
    210 : wave = 39010;
    211 : wave = 40812;
    212 : wave = 33206;
    213 : wave = 35055;
    214 : wave = 34873;
    215 : wave = 28579;
    216 : wave = 32810;
    217 : wave = 31921;
    218 : wave = 27043;
    219 : wave = 34173;
    220 : wave = 34013;
    221 : wave = 29505;
    222 : wave = 32176;
    223 : wave = 30340;
    224 : wave = 27798;
    225 : wave = 28514;
    226 : wave = 25611;
    227 : wave = 25143;
    228 : wave = 30453;
    229 : wave = 29187;
    230 : wave = 27885;
    231 : wave = 32789;
    232 : wave = 31278;
    233 : wave = 29762;
    234 : wave = 30963;
    235 : wave = 28218;
    236 : wave = 29039;
    237 : wave = 33914;
    238 : wave = 31776;
    239 : wave = 29895;
    240 : wave = 36074;
    241 : wave = 37779;
    242 : wave = 34297;
    243 : wave = 32363;
    244 : wave = 32868;
    245 : wave = 31655;
    246 : wave = 30534;
    247 : wave = 32966;
    248 : wave = 32882;
    249 : wave = 32107;
    250 : wave = 33273;
    251 : wave = 33828;
    252 : wave = 35940;
    253 : wave = 35441;
    254 : wave = 27813;
    255 : wave = 27384;
    256 : wave = 32394;
    257 : wave = 30998;
    258 : wave = 30418;
    259 : wave = 31904;
    260 : wave = 33195;
    261 : wave = 34742;
    262 : wave = 34532;
    263 : wave = 34234;
    264 : wave = 34352;
    265 : wave = 32052;
    266 : wave = 30351;
    267 : wave = 35118;
    268 : wave = 44261;
    269 : wave = 45396;
    270 : wave = 40045;
    271 : wave = 40255;
    272 : wave = 42611;
    273 : wave = 42864;
    274 : wave = 41763;
    275 : wave = 39076;
    276 : wave = 36459;
    277 : wave = 37359;
    278 : wave = 40917;
    279 : wave = 44541;
    280 : wave = 45869;
    281 : wave = 42881;
    282 : wave = 38455;
    283 : wave = 36712;
    284 : wave = 34600;
    285 : wave = 29296;
    286 : wave = 27964;
    287 : wave = 29884;
    288 : wave = 29217;
    289 : wave = 28121;
    290 : wave = 30035;
    291 : wave = 31811;
    292 : wave = 30744;
    293 : wave = 27465;
    294 : wave = 24395;
    295 : wave = 24018;
    296 : wave = 23439;
    297 : wave = 24511;
    298 : wave = 28196;
    299 : wave = 31307;
    300 : wave = 33010;
    301 : wave = 34419;
    302 : wave = 35166;
    303 : wave = 33770;
    304 : wave = 31513;
    305 : wave = 31323;
    306 : wave = 32685;
    307 : wave = 34045;
    308 : wave = 35324;
    309 : wave = 35421;
    310 : wave = 36933;
    311 : wave = 38343;
    312 : wave = 37516;
    313 : wave = 34710;
    314 : wave = 31289;
    315 : wave = 26997;
    316 : wave = 24227;
    317 : wave = 25480;
    318 : wave = 26080;
    319 : wave = 26458;
    320 : wave = 25375;
    321 : wave = 22738;
    322 : wave = 20101;
    323 : wave = 20018;
    324 : wave = 18670;
    325 : wave = 16247;
    326 : wave = 15589;
    327 : wave = 13864;
    328 : wave = 18453;
    329 : wave = 24018;
    330 : wave = 25794;
    331 : wave = 26945;
    332 : wave = 27877;
    333 : wave = 27444;
    334 : wave = 26968;
    335 : wave = 30433;
    336 : wave = 34443;
    337 : wave = 37426;
    338 : wave = 40155;
    339 : wave = 44371;
    340 : wave = 49200;
    341 : wave = 53062;
    342 : wave = 56173;
    343 : wave = 58058;
    344 : wave = 53431;
    345 : wave = 48042;
    346 : wave = 47662;
    347 : wave = 49816;
    348 : wave = 52790;
    349 : wave = 49192;
    350 : wave = 46606;
    351 : wave = 45159;
    352 : wave = 43264;
    353 : wave = 41744;
    354 : wave = 36079;
    355 : wave = 29617;
    356 : wave = 22589;
    357 : wave = 19882;
    358 : wave = 19326;
    359 : wave = 18428;
    360 : wave = 17750;
    361 : wave = 17849;
    362 : wave = 18955;
    363 : wave = 14962;
    364 : wave = 11520;
    365 : wave = 14758;
    366 : wave = 17301;
    367 : wave = 14697;
    368 : wave = 12779;
    369 : wave = 16238;
    370 : wave = 22538;
    371 : wave = 27247;
    372 : wave = 30464;
    373 : wave = 31726;
    374 : wave = 32783;
    375 : wave = 32104;
    376 : wave = 31790;
    377 : wave = 36824;
    378 : wave = 37490;
    379 : wave = 34533;
    380 : wave = 34129;
    381 : wave = 35043;
    382 : wave = 36523;
    383 : wave = 35981;
    384 : wave = 32214;
    385 : wave = 29496;
    386 : wave = 28599;
    387 : wave = 25827;
    388 : wave = 24044;
    389 : wave = 24023;
    390 : wave = 21778;
    391 : wave = 18817;
    392 : wave = 19021;
    393 : wave = 18225;
    394 : wave = 16618;
    395 : wave = 16545;
    396 : wave = 15531;
    397 : wave = 17387;
    398 : wave = 21026;
    399 : wave = 22082;
    400 : wave = 23135;
    401 : wave = 26068;
    402 : wave = 30068;
    403 : wave = 32017;
    404 : wave = 31443;
    405 : wave = 32449;
    406 : wave = 36740;
    407 : wave = 41835;
    408 : wave = 43696;
    409 : wave = 45036;
    410 : wave = 48751;
    411 : wave = 52626;
    412 : wave = 53387;
    413 : wave = 51156;
    414 : wave = 49150;
    415 : wave = 50584;
    416 : wave = 51690;
    417 : wave = 49322;
    418 : wave = 49996;
    419 : wave = 51998;
    420 : wave = 59846;
    421 : wave = 65536;
    422 : wave = 55584;
    423 : wave = 46104;
    424 : wave = 50686;
    425 : wave = 55514;
    426 : wave = 50624;
    427 : wave = 41088;
    428 : wave = 35119;
    429 : wave = 43907;
    430 : wave = 49682;
    431 : wave = 44581;
    432 : wave = 42347;
    433 : wave = 40049;
    434 : wave = 35820;
    435 : wave = 29992;
    436 : wave = 26818;
    437 : wave = 23977;
    438 : wave = 24000;
    439 : wave = 23966;
    440 : wave = 20463;
    441 : wave = 20249;
    442 : wave = 20666;
    443 : wave = 23509;
    444 : wave = 25740;
    445 : wave = 19012;
    446 : wave = 9382 ;
    447 : wave = 10176;
    448 : wave = 18148;
    449 : wave = 22543;
    450 : wave = 21530;
    451 : wave = 19496;
    452 : wave = 21020;
    453 : wave = 26425;
    454 : wave = 27835;
    455 : wave = 25059;
    456 : wave = 24316;
    457 : wave = 22650;
    458 : wave = 22500;
    459 : wave = 23486;
    460 : wave = 24899;
    461 : wave = 26522;
    462 : wave = 26353;
    463 : wave = 24575;
    464 : wave = 22312;
    465 : wave = 20956;
    466 : wave = 20674;
    467 : wave = 21687;
    468 : wave = 20997;
    469 : wave = 19941;
    470 : wave = 18733;
    471 : wave = 20289;
    472 : wave = 23204;
    473 : wave = 21968;
    474 : wave = 20190;
    475 : wave = 19207;
    476 : wave = 19496;
    477 : wave = 22779;
    478 : wave = 26640;
    479 : wave = 28927;
    480 : wave = 30702;
    481 : wave = 32377;
    482 : wave = 36007;
    483 : wave = 37892;
    484 : wave = 36724;
    485 : wave = 37626;
    486 : wave = 40200;
    487 : wave = 42875;
    488 : wave = 45321;
    489 : wave = 47964;
    490 : wave = 50173;
    491 : wave = 52343;
    492 : wave = 53935;
    493 : wave = 52294;
    494 : wave = 49353;
    495 : wave = 48228;
    496 : wave = 48428;
    497 : wave = 48620;
    498 : wave = 47082;
    499 : wave = 46412;
    500 : wave = 49336;
    501 : wave = 49865;
    502 : wave = 46330;
    503 : wave = 44036;
    504 : wave = 43086;
    505 : wave = 39370;
    506 : wave = 37850;
    507 : wave = 40476;
    508 : wave = 39781;
    509 : wave = 38406;
    510 : wave = 44905;
    511 : wave = 47578;
    512 : wave = 41127;
    513 : wave = 39802;
    514 : wave = 42831;
    515 : wave = 45541;
    516 : wave = 41213;
    517 : wave = 35346;
    518 : wave = 39608;
    519 : wave = 46354;
    520 : wave = 46179;
    521 : wave = 40928;
    522 : wave = 41358;
    523 : wave = 41183;
    524 : wave = 36267;
    525 : wave = 33146;
    526 : wave = 28933;
    527 : wave = 27168;
    528 : wave = 26464;
    529 : wave = 23338;
    530 : wave = 23144;
    531 : wave = 24984;
    532 : wave = 22331;
    533 : wave = 17059;
    534 : wave = 15826;
    535 : wave = 14208;
    536 : wave = 11959;
    537 : wave = 10896;
    538 : wave = 10501;
    539 : wave = 15312;
    540 : wave = 18240;
    541 : wave = 12422;
    542 : wave = 12348;
    543 : wave = 20793;
    544 : wave = 20210;
    545 : wave = 15184;
    546 : wave = 15184;
    547 : wave = 20475;
    548 : wave = 26792;
    549 : wave = 27441;
    550 : wave = 25726;
    551 : wave = 30096;
    552 : wave = 36428;
    553 : wave = 32179;
    554 : wave = 30110;
    555 : wave = 33302;
    556 : wave = 31294;
    557 : wave = 30323;
    558 : wave = 34048;
    559 : wave = 37203;
    560 : wave = 37231;
    561 : wave = 36061;
    562 : wave = 36729;
    563 : wave = 40399;
    564 : wave = 39054;
    565 : wave = 34988;
    566 : wave = 33529;
    567 : wave = 36419;
    568 : wave = 39004;
    569 : wave = 39280;
    570 : wave = 40786;
    571 : wave = 40463;
    572 : wave = 41445;
    573 : wave = 38825;
    574 : wave = 38180;
    575 : wave = 40864;
    576 : wave = 40045;
    577 : wave = 39682;
    578 : wave = 39938;
    579 : wave = 41690;
    580 : wave = 44551;
    581 : wave = 48658;
    582 : wave = 47891;
    583 : wave = 44915;
    584 : wave = 42382;
    585 : wave = 42903;
    586 : wave = 45549;
    587 : wave = 43853;
    588 : wave = 44850;
    589 : wave = 43420;
    590 : wave = 40818;
    591 : wave = 43577;
    592 : wave = 48054;
    593 : wave = 46241;
    594 : wave = 41230;
    595 : wave = 35397;
    596 : wave = 33111;
    597 : wave = 40229;
    598 : wave = 37104;
    599 : wave = 30186;
    600 : wave = 28250;
    601 : wave = 30226;
    602 : wave = 31628;
    603 : wave = 28701;
    604 : wave = 26620;
    605 : wave = 21284;
    606 : wave = 20269;
    607 : wave = 19841;
    608 : wave = 18730;
    609 : wave = 19779;
    610 : wave = 19560;
    611 : wave = 18458;
    612 : wave = 21549;
    613 : wave = 21534;
    614 : wave = 20204;
    615 : wave = 23637;
    616 : wave = 23674;
    617 : wave = 24533;
    618 : wave = 22204;
    619 : wave = 27314;
    620 : wave = 28370;
    621 : wave = 28643;
    622 : wave = 37545;
    623 : wave = 41883;
    624 : wave = 43962;
    625 : wave = 35006;
    626 : wave = 33367;
    627 : wave = 45182;
    628 : wave = 49278;
    629 : wave = 37991;
    630 : wave = 39506;
    631 : wave = 42568;
    632 : wave = 38333;
    633 : wave = 49766;
    634 : wave = 61128;
    635 : wave = 65495;
    636 : wave = 53596;
    637 : wave = 43739;
    638 : wave = 45301;
    639 : wave = 53854;
    640 : wave = 56333;
    641 : wave = 49877;
    642 : wave = 52369;
    643 : wave = 52468;
    644 : wave = 48330;
    645 : wave = 54623;
    646 : wave = 65536;
    647 : wave = 56852;
    648 : wave = 48294;
    649 : wave = 33760;
    650 : wave = 25495;
    651 : wave = 40707;
    652 : wave = 41690;
    653 : wave = 37289;
    654 : wave = 33312;
    655 : wave = 29046;
    656 : wave = 25285;
    657 : wave = 25759;
    658 : wave = 25836;
    659 : wave = 19113;
    660 : wave = 9461 ;
    661 : wave = 2281 ;
    662 : wave = 6056 ;
    663 : wave = 14836;
    664 : wave = 23411;
    665 : wave = 26472;
    666 : wave = 23869;
    667 : wave = 17890;
    668 : wave = 15248;
    669 : wave = 17710;
    670 : wave = 23887;
    671 : wave = 23675;
    672 : wave = 19924;
    673 : wave = 20458;
    674 : wave = 25164;
    675 : wave = 35937;
    676 : wave = 36996;
    677 : wave = 32855;
    678 : wave = 28982;
    679 : wave = 25332;
    680 : wave = 24079;
    681 : wave = 25332;
    682 : wave = 25762;
    683 : wave = 25230;
    684 : wave = 25785;
    685 : wave = 21472;
    686 : wave = 20629;
    687 : wave = 24249;
    688 : wave = 24331;
    689 : wave = 18951;
    690 : wave = 18577;
    691 : wave = 19836;
    692 : wave = 18034;
    693 : wave = 23487;
    694 : wave = 28660;
    695 : wave = 27908;
    696 : wave = 25901;
    697 : wave = 23944;
    698 : wave = 26773;
    699 : wave = 34324;
    700 : wave = 35050;
    701 : wave = 31755;
    702 : wave = 35652;
    703 : wave = 43727;
    704 : wave = 42932;
    705 : wave = 38409;
    706 : wave = 36660;
    707 : wave = 37379;
    708 : wave = 41993;
    709 : wave = 39480;
    710 : wave = 39099;
    711 : wave = 43898;
    712 : wave = 42984;
    713 : wave = 44674;
    714 : wave = 46907;
    715 : wave = 41526;
    716 : wave = 35093;
    717 : wave = 35101;
    718 : wave = 37591;
    719 : wave = 34901;
    720 : wave = 35186;
    721 : wave = 38456;
    722 : wave = 37803;
    723 : wave = 39521;
    724 : wave = 37699;
    725 : wave = 33750;
    726 : wave = 34797;
    727 : wave = 33493;
    728 : wave = 30332;
    729 : wave = 32142;
    730 : wave = 33499;
    731 : wave = 32539;
    732 : wave = 34434;
    733 : wave = 36170;
    734 : wave = 33374;
    735 : wave = 28622;
    736 : wave = 26780;
    737 : wave = 26934;
    738 : wave = 28250;
    739 : wave = 24278;
    740 : wave = 22918;
    741 : wave = 28298;
    742 : wave = 26472;
    743 : wave = 22384;
    744 : wave = 21490;
    745 : wave = 21377;
    746 : wave = 18092;
    747 : wave = 16169;
    748 : wave = 19900;
    749 : wave = 20413;
    750 : wave = 19482;
    751 : wave = 19081;
    752 : wave = 19024;
    753 : wave = 22569;
    754 : wave = 17602;
    755 : wave = 11506;
    756 : wave = 19038;
    757 : wave = 26023;
    758 : wave = 26377;
    759 : wave = 26492;
    760 : wave = 28570;
    761 : wave = 31295;
    762 : wave = 30416;
    763 : wave = 28022;
    764 : wave = 30050;
    765 : wave = 29296;
    766 : wave = 23988;
    767 : wave = 26116;
    768 : wave = 32525;
    769 : wave = 35772;
    770 : wave = 36471;
    771 : wave = 33657;
    772 : wave = 31100;
    773 : wave = 28359;
    774 : wave = 24760;
    775 : wave = 23107;
    776 : wave = 22204;
    777 : wave = 26918;
    778 : wave = 26019;
    779 : wave = 21502;
    780 : wave = 28219;
    781 : wave = 33384;
    782 : wave = 30781;
    783 : wave = 23835;
    784 : wave = 20809;
    785 : wave = 24185;
    786 : wave = 27226;
    787 : wave = 29162;
    788 : wave = 32879;
    789 : wave = 36506;
    790 : wave = 37760;
    791 : wave = 39591;
    792 : wave = 42364;
    793 : wave = 44833;
    794 : wave = 42289;
    795 : wave = 40170;
    796 : wave = 41929;
    797 : wave = 46130;
    798 : wave = 48020;
    799 : wave = 45108;
    800 : wave = 46568;
    801 : wave = 48306;
    802 : wave = 46185;
    803 : wave = 43521;
    804 : wave = 44139;
    805 : wave = 44430;
    806 : wave = 44718;
    807 : wave = 42732;
    808 : wave = 36880;
    809 : wave = 40618;
    810 : wave = 43582;
    811 : wave = 37619;
    812 : wave = 31666;
    813 : wave = 29196;
    814 : wave = 32940;
    815 : wave = 36616;
    816 : wave = 33395;
    817 : wave = 31098;
    818 : wave = 33747;
    819 : wave = 35946;
    820 : wave = 34751;
    821 : wave = 31436;
    822 : wave = 30949;
    823 : wave = 31861;
    824 : wave = 32348;
    825 : wave = 32206;
    826 : wave = 33242;
    827 : wave = 37524;
    828 : wave = 38540;
    829 : wave = 35211;
    830 : wave = 35269;
    831 : wave = 36608;
    832 : wave = 34622;
    833 : wave = 32640;
    834 : wave = 31202;
    835 : wave = 31054;
    836 : wave = 31513;
    837 : wave = 33520;
    838 : wave = 35591;
    839 : wave = 33671;
    840 : wave = 27371;
    841 : wave = 23866;
    842 : wave = 28672;
    843 : wave = 29437;
    844 : wave = 24919;
    845 : wave = 21255;
    846 : wave = 20225;
    847 : wave = 21896;
    848 : wave = 21820;
    849 : wave = 21685;
    850 : wave = 24739;
    851 : wave = 28228;
    852 : wave = 25978;
    853 : wave = 21057;
    854 : wave = 22035;
    855 : wave = 31091;
    856 : wave = 36019;
    857 : wave = 29315;
    858 : wave = 22697;
    859 : wave = 26989;
    860 : wave = 37031;
    861 : wave = 37882;
    862 : wave = 33625;
    863 : wave = 35313;
    864 : wave = 39234;
    865 : wave = 38973;
    866 : wave = 37486;
    867 : wave = 39659;
    868 : wave = 39317;
    869 : wave = 36856;
    870 : wave = 36799;
    871 : wave = 36538;
    872 : wave = 36018;
    873 : wave = 37167;
    874 : wave = 41299;
    875 : wave = 40786;
    876 : wave = 33615;
    877 : wave = 29927;
    878 : wave = 32070;
    879 : wave = 34030;
    880 : wave = 31503;
    881 : wave = 31922;
    882 : wave = 34526;
    883 : wave = 35464;
    884 : wave = 36878;
    885 : wave = 34939;
    886 : wave = 34152;
    887 : wave = 36074;
    888 : wave = 35882;
    889 : wave = 33175;
    890 : wave = 32804;
    891 : wave = 37205;
    892 : wave = 41624;
    893 : wave = 40699;
    894 : wave = 38456;
    895 : wave = 39680;
    896 : wave = 36129;
    897 : wave = 34428;
    898 : wave = 38261;
    899 : wave = 38784;
    900 : wave = 35545;
    901 : wave = 31370;
    902 : wave = 34590;
    903 : wave = 40696;
    904 : wave = 39270;
    905 : wave = 31692;
    906 : wave = 27743;
    907 : wave = 29505;
    908 : wave = 27873;
    909 : wave = 25231;
    910 : wave = 27590;
    911 : wave = 31442;
    912 : wave = 31343;
    913 : wave = 26422;
    914 : wave = 23724;
    915 : wave = 29583;
    916 : wave = 32009;
    917 : wave = 26516;
    918 : wave = 24139;
    919 : wave = 25683;
    920 : wave = 28869;
    921 : wave = 32148;
    922 : wave = 35063;
    923 : wave = 34066;
    924 : wave = 29956;
    925 : wave = 27593;
    926 : wave = 27929;
    927 : wave = 31492;
    928 : wave = 32797;
    929 : wave = 30677;
    930 : wave = 32055;
    931 : wave = 36701;
    932 : wave = 36634;
    933 : wave = 33627;
    934 : wave = 31813;
    935 : wave = 31753;
    936 : wave = 29881;
    937 : wave = 26737;
    938 : wave = 28549;
    939 : wave = 31929;
    940 : wave = 33555;
    941 : wave = 32482;
    942 : wave = 33813;
    943 : wave = 30744;
    944 : wave = 25660;
    945 : wave = 28507;
    946 : wave = 31398;
    947 : wave = 31449;
    948 : wave = 28733;
    949 : wave = 33720;
    950 : wave = 39549;
    951 : wave = 38987;
    952 : wave = 35775;
    953 : wave = 33134;
    954 : wave = 37208;
    955 : wave = 35482;
    956 : wave = 31941;
    957 : wave = 35282;
    958 : wave = 39547;
    959 : wave = 42079;
    960 : wave = 44828;
    961 : wave = 45304;
    962 : wave = 44139;
    963 : wave = 40547;
    964 : wave = 34947;
    965 : wave = 35047;
    966 : wave = 34164;
    967 : wave = 34474;
    968 : wave = 36798;
    969 : wave = 39512;
    970 : wave = 40538;
    971 : wave = 37480;
    972 : wave = 35119;
    973 : wave = 32878;
    974 : wave = 31100;
    975 : wave = 26878;
    976 : wave = 26593;
    977 : wave = 30096;
    978 : wave = 32742;
    979 : wave = 35302;
    980 : wave = 36349;
    981 : wave = 34211;
    982 : wave = 32098;
    983 : wave = 33303;
    984 : wave = 29840;
    985 : wave = 27015;
    986 : wave = 27508;
    987 : wave = 28950;
    988 : wave = 32777;
    989 : wave = 36593;
    990 : wave = 37159;
    991 : wave = 36169;
    992 : wave = 36274;
    993 : wave = 33392;
    994 : wave = 32208;
    995 : wave = 30162;
    996 : wave = 28472;
    997 : wave = 32299;
    998 : wave = 35662;
    999 : wave = 36569;
    1000: wave = 34928;
    1001: wave = 32962;
    1002: wave = 31784;
    1003: wave = 32107;
    1004: wave = 30519;
    1005: wave = 28456;
    1006: wave = 30769;
    1007: wave = 33728;
    1008: wave = 34960;
    1009: wave = 34336;
    1010: wave = 34530;
    1011: wave = 33578;
    1012: wave = 30984;
    1013: wave = 27546;
    1014: wave = 25155;
    1015: wave = 29745;
    1016: wave = 32574;
    1017: wave = 32522;
    1018: wave = 33927;
    1019: wave = 34101;
    1020: wave = 33474;
    1021: wave = 31526;
    1022: wave = 30676;
    1023: wave = 30485;
    1024: wave = 29078;
    1025: wave = 26611;
    1026: wave = 30940;
    1027: wave = 38418;
    1028: wave = 37994;
    1029: wave = 33578;
    1030: wave = 31893;
    1031: wave = 34202;
    1032: wave = 32708;
    1033: wave = 30229;
    1034: wave = 30673;
    1035: wave = 32089;
    1036: wave = 32141;
    1037: wave = 33903;
    1038: wave = 38479;
    1039: wave = 37954;
    1040: wave = 33651;
    1041: wave = 29603;
    1042: wave = 30950;
    1043: wave = 32984;
    1044: wave = 34461;
    1045: wave = 33840;
    1046: wave = 33189;
    1047: wave = 36268;
    1048: wave = 34857;
    1049: wave = 32978;
    1050: wave = 33384;
    1051: wave = 34606;
    1052: wave = 32542;
    1053: wave = 33306;
    1054: wave = 36148;
    1055: wave = 38145;
    1056: wave = 39566;
    1057: wave = 35610;
    1058: wave = 34039;
    1059: wave = 30964;
    1060: wave = 29707;
    1061: wave = 31977;
    1062: wave = 34875;
    1063: wave = 34594;
    1064: wave = 31365;
    1065: wave = 34066;
    1066: wave = 36189;
    1067: wave = 36799;
    1068: wave = 33868;
    1069: wave = 28544;
    1070: wave = 26637;
    1071: wave = 30036;
    1072: wave = 33352;
    1073: wave = 34521;
    1074: wave = 35975;
    1075: wave = 35104;
    1076: wave = 37725;
    1077: wave = 37722;
    1078: wave = 32772;
    1079: wave = 30805;
    1080: wave = 32017;
    1081: wave = 32447;
    1082: wave = 31460;
    1083: wave = 32975;
    1084: wave = 35609;
    1085: wave = 38871;
    1086: wave = 39710;
    1087: wave = 34373;
    1088: wave = 28254;
    1089: wave = 28240;
    1090: wave = 29092;
    1091: wave = 26911;
    1092: wave = 24572;
    1093: wave = 23886;
    1094: wave = 27029;
    1095: wave = 28952;
    1096: wave = 29022;
    1097: wave = 28767;
    1098: wave = 27676;
    1099: wave = 28004;
    1100: wave = 27206;
    1101: wave = 26081;
    1102: wave = 26457;
    1103: wave = 27970;
    1104: wave = 29818;
    1105: wave = 29501;
    1106: wave = 32293;
    1107: wave = 38156;
    1108: wave = 37745;
    1109: wave = 35182;
    1110: wave = 36558;
    1111: wave = 38124;
    1112: wave = 38526;
    1113: wave = 37516;
    1114: wave = 36691;
    1115: wave = 36476;
    1116: wave = 36280;
    1117: wave = 38166;
    1118: wave = 39784;
    1119: wave = 39233;
    1120: wave = 37046;
    1121: wave = 35821;
    1122: wave = 34387;
    1123: wave = 31890;
    1124: wave = 32237;
    1125: wave = 33012;
    1126: wave = 31613;
    1127: wave = 29772;
    1128: wave = 30427;
    1129: wave = 32011;
    1130: wave = 32922;
    1131: wave = 34111;
    1132: wave = 33038;
    1133: wave = 29582;
    1134: wave = 28591;
    1135: wave = 29913;
    1136: wave = 31434;
    1137: wave = 34065;
    1138: wave = 34707;
    1139: wave = 34085;
    1140: wave = 33932;
    1141: wave = 35643;
    1142: wave = 37522;
    1143: wave = 36895;
    1144: wave = 36549;
    1145: wave = 35899;
    1146: wave = 35914;
    1147: wave = 35299;
    1148: wave = 34849;
    1149: wave = 37783;
    1150: wave = 38023;
    1151: wave = 33567;
    1152: wave = 32987;
    1153: wave = 35356;
    1154: wave = 35716;
    1155: wave = 35557;
    1156: wave = 34324;
    1157: wave = 32833;
    1158: wave = 29942;
    1159: wave = 29116;
    1160: wave = 30229;
    1161: wave = 29344;
    1162: wave = 28955;
    1163: wave = 29255;
    1164: wave = 31285;
    1165: wave = 31883;
    1166: wave = 29917;
    1167: wave = 29837;
    1168: wave = 31961;
    1169: wave = 32453;
    1170: wave = 31550;
    1171: wave = 31262;
    1172: wave = 30130;
    1173: wave = 30775;
    1174: wave = 32742;
    1175: wave = 34049;
    1176: wave = 35638;
    1177: wave = 34317;
    1178: wave = 31434;
    1179: wave = 33357;
    1180: wave = 37182;
    1181: wave = 36622;
    1182: wave = 33514;
    1183: wave = 32792;
    1184: wave = 32902;
    1185: wave = 31800;
    1186: wave = 33265;
    1187: wave = 35519;
    1188: wave = 35137;
    1189: wave = 31622;
    1190: wave = 27723;
    1191: wave = 28463;
    1192: wave = 30709;
    1193: wave = 31774;
    1194: wave = 30650;
    1195: wave = 28472;
    1196: wave = 28367;
    1197: wave = 29435;
    1198: wave = 32261;
    1199: wave = 33248;
    1200: wave = 32666;
    1201: wave = 31517;
    1202: wave = 28507;
    1203: wave = 27517;
    1204: wave = 29272;
    1205: wave = 32261;
    1206: wave = 33604;
    1207: wave = 34237;
    1208: wave = 34837;
    1209: wave = 36955;
    1210: wave = 38716;
    1211: wave = 38175;
    1212: wave = 37416;
    1213: wave = 34878;
    1214: wave = 33767;
    1215: wave = 33544;
    1216: wave = 35870;
    1217: wave = 37896;
    1218: wave = 36918;
    1219: wave = 36199;
    1220: wave = 34693;
    1221: wave = 34858;
    1222: wave = 33921;
    1223: wave = 31597;
    1224: wave = 30891;
    1225: wave = 30999;
    1226: wave = 29089;
    1227: wave = 27255;
    1228: wave = 27085;
    1229: wave = 27767;
    1230: wave = 28715;
    1231: wave = 27281;
    1232: wave = 27142;
    1233: wave = 28520;
    1234: wave = 29937;
    1235: wave = 29377;
    1236: wave = 28622;
    1237: wave = 29785;
    1238: wave = 32160;
    1239: wave = 33459;
    1240: wave = 32110;
    1241: wave = 33168;
    1242: wave = 34733;
    1243: wave = 36868;
    1244: wave = 38488;
    1245: wave = 39210;
    1246: wave = 38949;
    1247: wave = 36445;
    1248: wave = 35760;
    1249: wave = 35855;
    1250: wave = 35636;
    1251: wave = 34942;
    1252: wave = 34846;
    1253: wave = 34695;
    1254: wave = 33248;
    1255: wave = 30595;
    1256: wave = 29061;
    1257: wave = 29437;
    1258: wave = 28619;
    1259: wave = 25746;
    1260: wave = 23440;
    1261: wave = 24743;
    1262: wave = 27076;
    1263: wave = 30097;
    1264: wave = 30641;
    1265: wave = 28041;
    1266: wave = 26673;
    1267: wave = 26312;
    1268: wave = 27082;
    1269: wave = 27905;
    1270: wave = 28648;
    1271: wave = 30975;
    1272: wave = 34149;
    1273: wave = 35772;
    1274: wave = 37341;
    1275: wave = 37792;
    1276: wave = 35299;
    1277: wave = 33560;
    1278: wave = 34056;
    1279: wave = 33808;
    1280: wave = 32902;
    1281: wave = 35969;
    1282: wave = 40019;
    1283: wave = 39489;
    1284: wave = 36322;
    1285: wave = 34103;
    1286: wave = 33712;
    1287: wave = 33815;
    1288: wave = 31129;
    1289: wave = 28015;
    1290: wave = 28952;
    1291: wave = 31492;
    1292: wave = 33024;
    1293: wave = 33590;
    1294: wave = 33540;
    1295: wave = 32830;
    1296: wave = 31262;
    1297: wave = 28620;
    1298: wave = 27603;
    1299: wave = 28361;
    1300: wave = 29151;
    1301: wave = 31652;
    1302: wave = 34565;
    1303: wave = 34559;
    1304: wave = 33032;
    1305: wave = 33453;
    1306: wave = 34259;
    1307: wave = 33930;
    1308: wave = 32597;
    1309: wave = 33020;
    1310: wave = 35879;
    1311: wave = 37724;
    1312: wave = 37463;
    1313: wave = 35293;
    1314: wave = 34832;
    1315: wave = 34753;
    1316: wave = 32244;
    1317: wave = 31980;
    1318: wave = 34429;
    1319: wave = 34303;
    1320: wave = 32557;
    1321: wave = 33343;
    1322: wave = 34863;
    1323: wave = 33767;
    1324: wave = 31256;
    1325: wave = 29858;
    1326: wave = 29121;
    1327: wave = 29747;
    1328: wave = 31123;
    1329: wave = 32237;
    1330: wave = 33747;
    1331: wave = 34706;
    1332: wave = 34854;
    1333: wave = 34124;
    1334: wave = 33697;
    1335: wave = 35070;
    1336: wave = 35087;
    1337: wave = 32882;
    1338: wave = 33285;
    1339: wave = 36088;
    1340: wave = 39219;
    1341: wave = 39663;
    1342: wave = 37173;
    1343: wave = 35685;
    1344: wave = 35527;
    1345: wave = 37013;
    1346: wave = 36422;
    1347: wave = 35075;
    1348: wave = 34455;
    1349: wave = 32785;
    1350: wave = 33227;
    1351: wave = 32971;
    1352: wave = 31700;
    1353: wave = 30320;
    1354: wave = 29753;
    1355: wave = 31896;
    1356: wave = 33203;
    1357: wave = 32881;
    1358: wave = 32315;
    1359: wave = 30593;
    1360: wave = 27778;
    1361: wave = 26440;
    1362: wave = 26000;
    1363: wave = 26094;
    1364: wave = 27401;
    1365: wave = 31816;
    1366: wave = 36235;
    1367: wave = 34458;
    1368: wave = 32823;
    1369: wave = 34951;
    1370: wave = 37109;
    1371: wave = 33993;
    1372: wave = 29057;
    1373: wave = 32168;
    1374: wave = 37649;
    1375: wave = 36286;
    1376: wave = 34242;
    1377: wave = 39144;
    1378: wave = 42070;
    1379: wave = 39738;
    1380: wave = 36700;
    1381: wave = 34686;
    1382: wave = 33410;
    1383: wave = 29711;
    1384: wave = 30285;
    1385: wave = 35119;
    1386: wave = 35881;
    1387: wave = 33097;
    1388: wave = 31619;
    1389: wave = 33917;
    1390: wave = 34858;
    1391: wave = 28497;
    1392: wave = 23472;
    1393: wave = 27656;
    1394: wave = 32101;
    1395: wave = 30294;
    1396: wave = 26289;
    1397: wave = 28396;
    1398: wave = 31774;
    1399: wave = 29476;
    1400: wave = 29559;
    1401: wave = 33265;
    1402: wave = 32713;
    1403: wave = 29672;
    1404: wave = 31492;
    1405: wave = 33448;
    1406: wave = 31791;
    1407: wave = 30326;
    1408: wave = 31889;
    1409: wave = 35215;
    1410: wave = 36607;
    1411: wave = 35195;
    1412: wave = 34237;
    1413: wave = 37390;
    1414: wave = 38580;
    1415: wave = 36451;
    1416: wave = 34434;
    1417: wave = 34606;
    1418: wave = 35856;
    1419: wave = 33494;
    1420: wave = 33003;
    1421: wave = 35154;
    1422: wave = 35859;
    1423: wave = 34594;
    1424: wave = 33636;
    1425: wave = 33219;
    1426: wave = 30093;
    1427: wave = 29283;
    1428: wave = 30184;
    1429: wave = 27789;
    1430: wave = 24691;
    1431: wave = 24249;
    1432: wave = 27189;
    1433: wave = 30761;
    1434: wave = 31762;
    1435: wave = 28283;
    1436: wave = 25611;
    1437: wave = 27018;
    1438: wave = 26631;
    1439: wave = 26452;
    1440: wave = 27238;
    1441: wave = 27894;
    1442: wave = 31427;
    1443: wave = 34762;
    1444: wave = 35792;
    1445: wave = 34780;
    1446: wave = 35699;
    1447: wave = 36614;
    1448: wave = 34266;
    1449: wave = 32684;
    1450: wave = 31475;
    1451: wave = 34785;
    1452: wave = 36351;
    1453: wave = 31387;
    1454: wave = 29812;
    1455: wave = 32052;
    1456: wave = 36622;
    1457: wave = 36029;
    1458: wave = 28912;
    1459: wave = 25350;
    1460: wave = 26477;
    1461: wave = 25926;
    1462: wave = 21960;
    1463: wave = 21844;
    1464: wave = 23703;
    1465: wave = 25697;
    1466: wave = 29299;
    1467: wave = 31648;
    1468: wave = 30668;
    1469: wave = 26959;
    1470: wave = 25778;
    1471: wave = 26429;
    1472: wave = 28564;
    1473: wave = 30998;
    1474: wave = 33732;
    1475: wave = 37495;
    1476: wave = 38722;
    1477: wave = 40048;
    1478: wave = 41178;
    1479: wave = 41789;
    1480: wave = 41778;
    1481: wave = 39524;
    1482: wave = 37635;
    1483: wave = 36933;
    1484: wave = 36389;
    1485: wave = 37214;
    1486: wave = 38356;
    1487: wave = 37054;
    1488: wave = 36169;
    1489: wave = 36459;
    1490: wave = 35447;
    1491: wave = 31427;
    1492: wave = 26000;
    1493: wave = 22888;
    1494: wave = 22737;
    1495: wave = 24707;
    1496: wave = 27716;
    1497: wave = 27278;
    1498: wave = 23873;
    1499: wave = 24778;
    1500: wave = 27757;
    1501: wave = 28034;
    1502: wave = 25041;
    1503: wave = 25724;
    1504: wave = 29751;
    1505: wave = 30517;
    1506: wave = 32133;
    1507: wave = 33824;
    1508: wave = 34878;
    1509: wave = 34411;
    1510: wave = 35154;
    1511: wave = 37951;
    1512: wave = 40017;
    1513: wave = 41696;
    1514: wave = 39666;
    1515: wave = 38186;
    1516: wave = 37905;
    1517: wave = 36941;
    1518: wave = 35772;
    1519: wave = 36579;
    1520: wave = 37727;
    1521: wave = 33404;
    1522: wave = 28865;
    1523: wave = 30497;
    1524: wave = 34956;
    1525: wave = 31423;
    1526: wave = 25273;
    1527: wave = 25256;
    1528: wave = 26951;
    1529: wave = 27088;
    1530: wave = 24285;
    1531: wave = 23556;
    1532: wave = 25991;
    1533: wave = 27822;
    1534: wave = 28582;
    1535: wave = 28759;
    1536: wave = 30044;
    1537: wave = 30809;
    1538: wave = 29983;
    1539: wave = 30851;
    1540: wave = 33709;
    1541: wave = 36825;
    1542: wave = 37573;
    1543: wave = 38778;
    1544: wave = 43530;
    1545: wave = 43597;
    1546: wave = 38027;
    1547: wave = 37071;
    1548: wave = 41920;
    1549: wave = 42684;
    1550: wave = 40884;
    1551: wave = 39729;
    1552: wave = 38772;
    1553: wave = 40486;
    1554: wave = 39964;
    1555: wave = 37017;
    1556: wave = 32989;
    1557: wave = 33001;
    1558: wave = 33773;
    1559: wave = 27876;
    1560: wave = 25024;
    1561: wave = 27046;
    1562: wave = 28709;
    1563: wave = 28523;
    1564: wave = 27571;
    1565: wave = 26626;
    1566: wave = 25038;
    1567: wave = 21977;
    1568: wave = 20576;
    1569: wave = 21781;
    1570: wave = 21310;
    1571: wave = 22929;
    1572: wave = 26145;
    1573: wave = 29153;
    1574: wave = 31750;
    1575: wave = 31565;
    1576: wave = 31573;
    1577: wave = 31964;
    1578: wave = 32073;
    1579: wave = 30653;
    1580: wave = 28836;
    1581: wave = 31500;
    1582: wave = 35516;
    1583: wave = 37966;
    1584: wave = 39372;
    1585: wave = 40385;
    1586: wave = 40969;
    1587: wave = 39730;
    1588: wave = 38391;
    1589: wave = 35911;
    1590: wave = 33078;
    1591: wave = 32449;
    1592: wave = 33148;
    1593: wave = 35456;
    1594: wave = 38464;
    1595: wave = 37709;
    1596: wave = 35098;
    1597: wave = 34202;
    1598: wave = 30552;
    1599: wave = 28179;
    1600: wave = 28791;
    1601: wave = 27360;
    1602: wave = 24804;
    1603: wave = 25402;
    1604: wave = 30230;
    1605: wave = 35343;
    1606: wave = 37522;
    1607: wave = 35641;
    1608: wave = 35813;
    1609: wave = 34307;
    1610: wave = 29681;
    1611: wave = 29481;
    1612: wave = 31890;
    1613: wave = 33668;
    1614: wave = 36041;
    1615: wave = 41285;
    1616: wave = 42053;
    1617: wave = 40319;
    1618: wave = 39431;
    1619: wave = 39396;
    1620: wave = 39541;
    1621: wave = 35731;
    1622: wave = 36291;
    1623: wave = 38148;
    1624: wave = 36744;
    1625: wave = 35939;
    1626: wave = 35856;
    1627: wave = 35787;
    1628: wave = 35881;
    1629: wave = 34999;
    1630: wave = 32505;
    1631: wave = 31993;
    1632: wave = 30799;
    1633: wave = 31114;
    1634: wave = 31817;
    1635: wave = 29171;
    1636: wave = 28547;
    1637: wave = 30052;
    1638: wave = 32943;
    1639: wave = 34951;
    1640: wave = 31182;
    1641: wave = 26371;
    1642: wave = 29187;
    1643: wave = 34255;
    1644: wave = 34773;
    1645: wave = 32669;
    1646: wave = 31121;
    1647: wave = 30731;
    1648: wave = 28186;
    1649: wave = 27020;
    1650: wave = 30879;
    1651: wave = 35986;
    1652: wave = 38108;
    1653: wave = 36648;
    1654: wave = 34634;
    1655: wave = 33108;
    1656: wave = 31335;
    1657: wave = 29725;
    1658: wave = 28898;
    1659: wave = 28335;
    1660: wave = 28298;
    1661: wave = 31230;
    1662: wave = 35043;
    1663: wave = 34640;
    1664: wave = 31570;
    1665: wave = 28881;
    1666: wave = 29031;
    1667: wave = 29730;
    1668: wave = 26228;
    1669: wave = 23947;
    1670: wave = 25433;
    1671: wave = 26577;
    1672: wave = 26289;
    1673: wave = 27903;
    1674: wave = 31300;
    1675: wave = 33103;
    1676: wave = 33029;
    1677: wave = 30268;
    1678: wave = 30149;
    1679: wave = 31948;
    1680: wave = 32763;
    1681: wave = 37576;
    1682: wave = 42649;
    1683: wave = 43443;
    1684: wave = 41835;
    1685: wave = 42349;
    1686: wave = 43232;
    1687: wave = 41928;
    1688: wave = 41632;
    1689: wave = 43284;
    1690: wave = 46162;
    1691: wave = 45555;
    1692: wave = 40713;
    1693: wave = 38883;
    1694: wave = 40492;
    1695: wave = 37782;
    1696: wave = 34124;
    1697: wave = 32974;
    1698: wave = 30912;
    1699: wave = 30308;
    1700: wave = 30604;
    1701: wave = 32279;
    1702: wave = 33100;
    1703: wave = 30606;
    1704: wave = 28395;
    1705: wave = 26986;
    1706: wave = 25570;
    1707: wave = 23992;
    1708: wave = 22891;
    1709: wave = 25914;
    1710: wave = 31863;
    1711: wave = 33166;
    1712: wave = 33799;
    1713: wave = 34068;
    1714: wave = 32546;
    1715: wave = 32646;
    1716: wave = 31672;
    1717: wave = 31927;
    1718: wave = 31192;
    1719: wave = 30566;
    1720: wave = 32778;
    1721: wave = 37129;
    1722: wave = 40127;
    1723: wave = 38731;
    1724: wave = 38581;
    1725: wave = 36398;
    1726: wave = 33325;
    1727: wave = 30409;
    1728: wave = 28532;
    1729: wave = 30749;
    1730: wave = 31004;
    1731: wave = 30699;
    1732: wave = 33277;
    1733: wave = 37214;
    1734: wave = 37159;
    1735: wave = 34091;
    1736: wave = 30361;
    1737: wave = 26400;
    1738: wave = 25027;
    1739: wave = 25633;
    1740: wave = 26655;
    1741: wave = 26625;
    1742: wave = 28941;
    1743: wave = 30863;
    1744: wave = 31642;
    1745: wave = 33462;
    1746: wave = 32978;
    1747: wave = 31835;
    1748: wave = 32276;
    1749: wave = 32917;
    1750: wave = 31303;
    1751: wave = 31095;
    1752: wave = 33854;
    1753: wave = 40646;
    1754: wave = 46321;
    1755: wave = 44491;
    1756: wave = 42572;
    1757: wave = 40275;
    1758: wave = 38043;
    1759: wave = 39050;
    1760: wave = 39285;
    1761: wave = 38842;
    1762: wave = 38598;
    1763: wave = 38775;
    1764: wave = 41615;
    1765: wave = 43333;
    1766: wave = 41098;
    1767: wave = 37916;
    1768: wave = 34556;
    1769: wave = 33412;
    1770: wave = 32966;
    1771: wave = 32489;
    1772: wave = 34065;
    1773: wave = 35083;
    1774: wave = 36488;
    1775: wave = 38540;
    1776: wave = 39869;
    1777: wave = 41967;
    1778: wave = 42112;
    1779: wave = 39694;
    1780: wave = 38854;
    1781: wave = 38449;
    1782: wave = 40202;
    1783: wave = 45309;
    1784: wave = 48155;
    1785: wave = 46505;
    1786: wave = 41764;
    1787: wave = 37562;
    1788: wave = 37957;
    1789: wave = 39654;
    1790: wave = 35168;
    1791: wave = 27862;
    1792: wave = 25480;
    1793: wave = 27268;
    1794: wave = 29283;
    1795: wave = 28091;
    1796: wave = 21936;
    1797: wave = 17018;
    1798: wave = 17546;
    1799: wave = 16169;
    1800: wave = 11729;
    1801: wave = 11798;
    1802: wave = 15431;
    1803: wave = 17141;
    1804: wave = 17489;
    1805: wave = 16914;
    1806: wave = 19203;
    1807: wave = 23951;
    1808: wave = 23606;
    1809: wave = 21284;
    1810: wave = 21000;
    1811: wave = 23564;
    1812: wave = 29475;
    1813: wave = 34422;
    1814: wave = 34388;
    1815: wave = 32624;
    1816: wave = 32106;
    1817: wave = 32885;
    1818: wave = 35691;
    1819: wave = 34298;
    1820: wave = 29724;
    1821: wave = 29441;
    1822: wave = 31108;
    1823: wave = 30047;
    1824: wave = 27766;
    1825: wave = 28771;
    1826: wave = 31094;
    1827: wave = 30715;
    1828: wave = 27909;
    1829: wave = 25247;
    1830: wave = 25608;
    1831: wave = 27503;
    1832: wave = 27960;
    1833: wave = 26724;
    1834: wave = 26341;
    1835: wave = 27914;
    1836: wave = 29083;
    1837: wave = 31106;
    1838: wave = 31985;
    1839: wave = 32974;
    1840: wave = 37348;
    1841: wave = 39549;
    1842: wave = 40158;
    1843: wave = 38603;
    1844: wave = 36560;
    1845: wave = 38771;
    1846: wave = 41130;
    1847: wave = 41954;
    1848: wave = 42597;
    1849: wave = 43710;
    1850: wave = 44003;
    1851: wave = 42309;
    1852: wave = 40135;
    1853: wave = 38406;
    1854: wave = 36528;
    1855: wave = 35290;
    1856: wave = 33477;
    1857: wave = 31239;
    1858: wave = 31079;
    1859: wave = 31454;
    1860: wave = 31584;
    1861: wave = 30632;
    1862: wave = 29287;
    1863: wave = 27062;
    1864: wave = 24104;
    1865: wave = 22753;
    1866: wave = 22703;
    1867: wave = 23631;
    1868: wave = 24389;
    1869: wave = 26368;
    1870: wave = 28793;
    1871: wave = 29255;
    1872: wave = 28959;
    1873: wave = 29252;
    1874: wave = 30320;
    1875: wave = 31387;
    1876: wave = 31535;
    1877: wave = 31469;
    1878: wave = 33102;
    1879: wave = 33598;
    1880: wave = 32537;
    1881: wave = 33067;
    1882: wave = 33250;
    1883: wave = 31762;
    1884: wave = 30203;
    1885: wave = 29150;
    1886: wave = 28796;
    1887: wave = 28898;
    1888: wave = 28536;
    1889: wave = 28054;
    1890: wave = 27984;
    1891: wave = 27612;
    1892: wave = 26550;
    1893: wave = 26251;
    1894: wave = 26461;
    1895: wave = 26368;
    1896: wave = 26626;
    1897: wave = 27420;
    1898: wave = 28884;
    1899: wave = 29882;
    1900: wave = 30372;
    1901: wave = 31105;
    1902: wave = 32415;
    1903: wave = 33905;
    1904: wave = 34548;
    1905: wave = 35494;
    1906: wave = 36431;
    1907: wave = 36944;
    1908: wave = 38087;
    1909: wave = 38887;
    1910: wave = 39857;
    1911: wave = 40803;
    1912: wave = 40753;
    1913: wave = 40138;
    1914: wave = 38883;
    1915: wave = 38624;
    1916: wave = 37947;
    1917: wave = 36840;
    1918: wave = 36404;
    1919: wave = 35801;
    1920: wave = 36412;
    1921: wave = 36814;
    1922: wave = 37519;
    1923: wave = 38127;
    1924: wave = 36996;
    1925: wave = 35473;
    1926: wave = 34591;
    1927: wave = 34146;
    1928: wave = 33116;
    1929: wave = 32807;
    1930: wave = 33271;
    1931: wave = 34759;
    1932: wave = 36592;
    1933: wave = 38476;
    1934: wave = 40188;
    1935: wave = 39625;
    1936: wave = 38352;
    1937: wave = 37530;
    1938: wave = 37524;
    1939: wave = 37960;
    1940: wave = 38458;
    1941: wave = 38392;
    1942: wave = 38421;
    1943: wave = 39274;
    1944: wave = 39411;
    1945: wave = 39721;
    1946: wave = 39334;
    1947: wave = 37971;
    1948: wave = 36288;
    1949: wave = 34233;
    1950: wave = 33195;
    1951: wave = 33343;
    1952: wave = 33325;
    1953: wave = 32865;
    1954: wave = 32865;
    1955: wave = 32218;
    1956: wave = 31620;
    1957: wave = 31051;
    1958: wave = 30017;
    1959: wave = 29283;
    1960: wave = 27517;
    1961: wave = 26947;
    1962: wave = 27426;
    1963: wave = 27305;
    1964: wave = 28605;
    1965: wave = 30216;
    1966: wave = 31436;
    1967: wave = 32301;
    1968: wave = 32720;
    1969: wave = 32513;
    1970: wave = 31469;
    1971: wave = 31330;
    1972: wave = 31648;
    1973: wave = 31834;
    1974: wave = 32124;
    1975: wave = 33221;
    1976: wave = 34832;
    1977: wave = 35700;
    1978: wave = 36387;
    1979: wave = 36300;
    1980: wave = 35673;
    1981: wave = 34967;
    1982: wave = 34136;
    1983: wave = 33682;
    1984: wave = 33782;
    1985: wave = 34359;
    1986: wave = 35302;
    1987: wave = 36393;
    1988: wave = 36712;
    1989: wave = 36581;
    1990: wave = 35913;
    1991: wave = 34686;
    1992: wave = 33262;
    1993: wave = 32046;
    1994: wave = 31616;
    1995: wave = 32327;
    1996: wave = 34106;
    1997: wave = 35171;
    1998: wave = 35874;
    1999: wave = 35919;
    2000: wave = 35206;
    2001: wave = 35502;
    2002: wave = 35339;
    2003: wave = 34675;
    2004: wave = 34861;
    2005: wave = 34815;
    2006: wave = 34780;
    2007: wave = 36157;
    2008: wave = 37626;
    2009: wave = 38212;
    2010: wave = 38229;
    2011: wave = 37748;
    2012: wave = 37539;
    2013: wave = 36965;
    2014: wave = 36151;
    2015: wave = 36145;
    2016: wave = 35845;
    2017: wave = 35119;
    2018: wave = 34921;
    2019: wave = 34838;
    2020: wave = 34396;
    2021: wave = 33990;
    2022: wave = 33491;
    2023: wave = 33024;
    2024: wave = 33116;
    2025: wave = 32308;
    2026: wave = 31228;
    2027: wave = 31126;
    2028: wave = 30552;
    2029: wave = 30030;
    2030: wave = 29959;
    2031: wave = 30499;
    2032: wave = 31243;
    2033: wave = 31181;
    2034: wave = 30995;
    2035: wave = 30297;
    2036: wave = 29985;
    2037: wave = 29840;
    2038: wave = 29217;
    2039: wave = 29174;
    2040: wave = 29202;
    2041: wave = 29754;
    2042: wave = 30316;
    2043: wave = 30728;
    2044: wave = 31155;
    2045: wave = 31031;
    2046: wave = 30807;
    2047: wave = 30226;
    2048: wave = 29888;
    2049: wave = 29830;
    2050: wave = 30091;
    2051: wave = 30554;
    2052: wave = 30905;
    2053: wave = 31433;
    2054: wave = 31611;
    2055: wave = 31546;
    2056: wave = 31175;
    2057: wave = 30714;
    2058: wave = 30685;
    2059: wave = 31196;
    2060: wave = 31845;
    2061: wave = 32618;
    2062: wave = 33232;
    2063: wave = 33366;
    2064: wave = 33558; 
    default	:wave =16'h7374;
endcase
end

endmodule