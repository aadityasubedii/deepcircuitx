module coeffs31(
  input wire [3:0] select,
  input wire [4:0] index,
  output reg signed [9:0] coeff
);