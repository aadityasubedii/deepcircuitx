    always @(posedge dqs_odd[13]) dqs_odd_receiver(13);