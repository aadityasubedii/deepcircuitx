        always @* begin
            reset_out = reset_out_pre;
            reset_req = reset_req_pre;
        end