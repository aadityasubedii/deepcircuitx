always @ ( posedge `U_SYSTEM.clk )
    clk_count <= clk_count + 1'd1;
