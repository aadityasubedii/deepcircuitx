    always @(negedge dqs_in[25]) dqs_pos_timing_check(25);