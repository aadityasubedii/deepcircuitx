    always @(posedge clk) sync_0 <= i_btn;