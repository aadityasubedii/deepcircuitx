always @(posedge CLOCK_50) blink_cnt++;
