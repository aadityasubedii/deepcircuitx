always @ (wr_en or Reset or Start)
begin