    always @(addr_in[13]) cmd_addr_timing_check(20);