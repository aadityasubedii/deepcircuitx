`endif 
endmodule